module xls_conv_top(
  input wire clk,
  input wire [255:0] signal,
  input wire [255:0] kernel,
  input wire [255:0] output,
  output wire [255:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] smul32b_16b_x_16b (input reg [15:0] lhs, input reg [15:0] rhs);
    reg signed [15:0] signed_lhs;
    reg signed [15:0] signed_rhs;
    reg signed [31:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul32b_16b_x_16b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [46:0] smul47b_16b_x_31b (input reg [15:0] lhs, input reg [30:0] rhs);
    reg signed [15:0] signed_lhs;
    reg signed [30:0] signed_rhs;
    reg signed [46:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul47b_16b_x_31b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [47:0] smul48b_16b_x_32b (input reg [15:0] lhs, input reg [31:0] rhs);
    reg signed [15:0] signed_lhs;
    reg signed [31:0] signed_rhs;
    reg signed [47:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul48b_16b_x_32b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [15:0] smul16b_16b_x_16b (input reg [15:0] lhs, input reg [15:0] rhs);
    reg signed [15:0] signed_lhs;
    reg signed [15:0] signed_rhs;
    reg signed [15:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul16b_16b_x_16b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [48:0] smul49b_16b_x_33b (input reg [15:0] lhs, input reg [32:0] rhs);
    reg signed [15:0] signed_lhs;
    reg signed [32:0] signed_rhs;
    reg signed [48:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul49b_16b_x_33b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  function automatic [31:0] sdiv_32b (input reg [31:0] lhs, input reg [31:0] rhs);
    begin
      sdiv_32b = rhs == 32'h0000_0000 ? (lhs[31] ? 32'h8000_0000 : 32'h7fff_ffff) : (lhs == 32'h8000_0000 && rhs == 32'hffff_ffff ? 32'h8000_0000 : $unsigned($signed(lhs) / $signed(rhs)));
    end
  endfunction
  wire [15:0] signal_unflattened[16];
  assign signal_unflattened[0] = signal[15:0];
  assign signal_unflattened[1] = signal[31:16];
  assign signal_unflattened[2] = signal[47:32];
  assign signal_unflattened[3] = signal[63:48];
  assign signal_unflattened[4] = signal[79:64];
  assign signal_unflattened[5] = signal[95:80];
  assign signal_unflattened[6] = signal[111:96];
  assign signal_unflattened[7] = signal[127:112];
  assign signal_unflattened[8] = signal[143:128];
  assign signal_unflattened[9] = signal[159:144];
  assign signal_unflattened[10] = signal[175:160];
  assign signal_unflattened[11] = signal[191:176];
  assign signal_unflattened[12] = signal[207:192];
  assign signal_unflattened[13] = signal[223:208];
  assign signal_unflattened[14] = signal[239:224];
  assign signal_unflattened[15] = signal[255:240];
  wire [15:0] kernel_unflattened[16];
  assign kernel_unflattened[0] = kernel[15:0];
  assign kernel_unflattened[1] = kernel[31:16];
  assign kernel_unflattened[2] = kernel[47:32];
  assign kernel_unflattened[3] = kernel[63:48];
  assign kernel_unflattened[4] = kernel[79:64];
  assign kernel_unflattened[5] = kernel[95:80];
  assign kernel_unflattened[6] = kernel[111:96];
  assign kernel_unflattened[7] = kernel[127:112];
  assign kernel_unflattened[8] = kernel[143:128];
  assign kernel_unflattened[9] = kernel[159:144];
  assign kernel_unflattened[10] = kernel[175:160];
  assign kernel_unflattened[11] = kernel[191:176];
  assign kernel_unflattened[12] = kernel[207:192];
  assign kernel_unflattened[13] = kernel[223:208];
  assign kernel_unflattened[14] = kernel[239:224];
  assign kernel_unflattened[15] = kernel[255:240];
  wire [15:0] output_unflattened[16];
  assign output_unflattened[0] = output[15:0];
  assign output_unflattened[1] = output[31:16];
  assign output_unflattened[2] = output[47:32];
  assign output_unflattened[3] = output[63:48];
  assign output_unflattened[4] = output[79:64];
  assign output_unflattened[5] = output[95:80];
  assign output_unflattened[6] = output[111:96];
  assign output_unflattened[7] = output[127:112];
  assign output_unflattened[8] = output[143:128];
  assign output_unflattened[9] = output[159:144];
  assign output_unflattened[10] = output[175:160];
  assign output_unflattened[11] = output[191:176];
  assign output_unflattened[12] = output[207:192];
  assign output_unflattened[13] = output[223:208];
  assign output_unflattened[14] = output[239:224];
  assign output_unflattened[15] = output[255:240];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [15:0] p0_signal[16];
  reg [15:0] p0_kernel[16];
  always_ff @ (posedge clk) begin
    p0_signal <= signal_unflattened;
    p0_kernel <= kernel_unflattened;
  end

  // ===== Pipe stage 1:
  wire [15:0] p1_array_index_36119_comb;
  wire [15:0] p1_array_index_36120_comb;
  wire [15:0] p1_array_index_36121_comb;
  wire [15:0] p1_array_index_36122_comb;
  wire [15:0] p1_array_index_36123_comb;
  wire [15:0] p1_array_index_36124_comb;
  wire [15:0] p1_array_index_36125_comb;
  wire [15:0] p1_array_index_36126_comb;
  wire [15:0] p1_array_index_36127_comb;
  wire [15:0] p1_array_index_36128_comb;
  wire [15:0] p1_array_index_36129_comb;
  wire [15:0] p1_array_index_36130_comb;
  wire [15:0] p1_array_index_36131_comb;
  wire [15:0] p1_array_index_36132_comb;
  wire [15:0] p1_array_index_36133_comb;
  wire [15:0] p1_array_index_36134_comb;
  wire [15:0] p1_array_index_36135_comb;
  wire [15:0] p1_array_index_36136_comb;
  wire [15:0] p1_array_index_36137_comb;
  wire [15:0] p1_array_index_36138_comb;
  wire [15:0] p1_array_index_36139_comb;
  wire [15:0] p1_array_index_36140_comb;
  wire [15:0] p1_array_index_36141_comb;
  wire [15:0] p1_array_index_36142_comb;
  wire [15:0] p1_array_index_36143_comb;
  wire [15:0] p1_array_index_36144_comb;
  wire [15:0] p1_array_index_36145_comb;
  wire [15:0] p1_array_index_36146_comb;
  wire [15:0] p1_array_index_36148_comb;
  wire [15:0] p1_array_index_36149_comb;
  wire [31:0] p1_smul_36151_comb;
  wire [31:0] p1_smul_36152_comb;
  wire [31:0] p1_smul_36153_comb;
  wire [31:0] p1_smul_36154_comb;
  wire [31:0] p1_smul_36155_comb;
  wire [31:0] p1_smul_36156_comb;
  wire [31:0] p1_smul_36157_comb;
  wire [31:0] p1_smul_36158_comb;
  wire [31:0] p1_smul_36159_comb;
  wire [31:0] p1_smul_36160_comb;
  wire [31:0] p1_smul_36161_comb;
  wire [31:0] p1_smul_36162_comb;
  wire [31:0] p1_smul_36163_comb;
  wire [31:0] p1_smul_36164_comb;
  wire [31:0] p1_smul_36165_comb;
  wire [31:0] p1_smul_36166_comb;
  wire [31:0] p1_smul_36167_comb;
  wire [31:0] p1_smul_36168_comb;
  wire [31:0] p1_smul_36169_comb;
  wire [31:0] p1_smul_36170_comb;
  wire [31:0] p1_smul_36171_comb;
  wire [31:0] p1_smul_36172_comb;
  wire [31:0] p1_smul_36173_comb;
  wire [31:0] p1_smul_36174_comb;
  wire [31:0] p1_smul_36175_comb;
  wire [31:0] p1_smul_36176_comb;
  wire [31:0] p1_smul_36177_comb;
  wire [31:0] p1_smul_36178_comb;
  wire [31:0] p1_smul_36179_comb;
  wire [31:0] p1_smul_36180_comb;
  wire [31:0] p1_smul_36181_comb;
  wire [31:0] p1_smul_36182_comb;
  wire [31:0] p1_smul_36183_comb;
  wire [31:0] p1_smul_36184_comb;
  wire [31:0] p1_smul_36185_comb;
  wire [31:0] p1_smul_36186_comb;
  wire [31:0] p1_smul_36187_comb;
  wire [31:0] p1_smul_36188_comb;
  wire [31:0] p1_smul_36189_comb;
  wire [31:0] p1_smul_36190_comb;
  wire [31:0] p1_smul_36191_comb;
  wire [31:0] p1_smul_36192_comb;
  wire [31:0] p1_smul_36193_comb;
  wire [31:0] p1_smul_36194_comb;
  wire [31:0] p1_smul_36195_comb;
  wire [31:0] p1_smul_36196_comb;
  wire [31:0] p1_smul_36197_comb;
  wire [31:0] p1_smul_36198_comb;
  wire [31:0] p1_smul_36199_comb;
  wire [31:0] p1_smul_36200_comb;
  wire [31:0] p1_smul_36201_comb;
  wire [31:0] p1_smul_36202_comb;
  wire [31:0] p1_smul_36203_comb;
  wire [31:0] p1_smul_36204_comb;
  wire [31:0] p1_smul_36205_comb;
  wire [31:0] p1_smul_36206_comb;
  wire [31:0] p1_smul_36207_comb;
  wire [31:0] p1_smul_36208_comb;
  wire [31:0] p1_smul_36209_comb;
  wire [31:0] p1_smul_36210_comb;
  wire [31:0] p1_smul_36211_comb;
  wire [31:0] p1_smul_36212_comb;
  wire [31:0] p1_smul_36213_comb;
  wire [31:0] p1_smul_36214_comb;
  wire [31:0] p1_smul_36215_comb;
  wire [31:0] p1_smul_36216_comb;
  wire [31:0] p1_smul_36217_comb;
  wire [31:0] p1_smul_36218_comb;
  wire [31:0] p1_smul_36219_comb;
  wire [31:0] p1_smul_36220_comb;
  wire [31:0] p1_smul_36221_comb;
  wire [31:0] p1_smul_36222_comb;
  wire [31:0] p1_smul_36223_comb;
  wire [31:0] p1_smul_36224_comb;
  wire [31:0] p1_smul_36225_comb;
  wire [31:0] p1_smul_36226_comb;
  wire [31:0] p1_smul_36227_comb;
  wire [31:0] p1_smul_36228_comb;
  wire [31:0] p1_smul_36229_comb;
  wire [31:0] p1_smul_36230_comb;
  wire [31:0] p1_smul_36231_comb;
  wire [31:0] p1_smul_36232_comb;
  wire [31:0] p1_smul_36233_comb;
  wire [31:0] p1_smul_36234_comb;
  wire [31:0] p1_smul_36235_comb;
  wire [31:0] p1_smul_36236_comb;
  wire [31:0] p1_smul_36237_comb;
  wire [31:0] p1_smul_36238_comb;
  wire [31:0] p1_smul_36239_comb;
  wire [31:0] p1_smul_36240_comb;
  wire [31:0] p1_smul_36241_comb;
  wire [31:0] p1_smul_36242_comb;
  wire [31:0] p1_smul_36245_comb;
  wire [31:0] p1_smul_36246_comb;
  wire [31:0] p1_smul_36247_comb;
  wire [31:0] p1_smul_36248_comb;
  wire [31:0] p1_smul_36249_comb;
  wire [31:0] p1_smul_36250_comb;
  wire [31:0] p1_smul_36251_comb;
  wire [31:0] p1_smul_36256_comb;
  wire [31:0] p1_smul_36257_comb;
  wire [31:0] p1_smul_36258_comb;
  wire [31:0] p1_smul_36259_comb;
  wire [31:0] p1_smul_36260_comb;
  wire [31:0] p1_smul_36261_comb;
  wire [31:0] p1_smul_36268_comb;
  wire [31:0] p1_smul_36269_comb;
  wire [31:0] p1_smul_36270_comb;
  wire [31:0] p1_smul_36271_comb;
  wire [31:0] p1_smul_36272_comb;
  wire [31:0] p1_smul_36281_comb;
  wire [31:0] p1_smul_36282_comb;
  wire [31:0] p1_smul_36283_comb;
  wire [31:0] p1_smul_36284_comb;
  wire [31:0] p1_smul_36295_comb;
  wire [31:0] p1_smul_36296_comb;
  wire [31:0] p1_smul_36297_comb;
  wire [31:0] p1_smul_36310_comb;
  wire [31:0] p1_smul_36311_comb;
  wire [31:0] p1_smul_36326_comb;
  wire [31:0] p1_smul_36343_comb;
  wire [31:0] p1_smul_36344_comb;
  wire [31:0] p1_smul_36345_comb;
  wire [31:0] p1_smul_36346_comb;
  wire [31:0] p1_smul_36347_comb;
  wire [31:0] p1_smul_36348_comb;
  wire [31:0] p1_smul_36351_comb;
  wire [31:0] p1_smul_36352_comb;
  wire [31:0] p1_smul_36353_comb;
  wire [31:0] p1_smul_36358_comb;
  wire [31:0] p1_smul_36359_comb;
  wire [31:0] p1_smul_36366_comb;
  wire [15:0] p1_add_36375_comb;
  wire [15:0] p1_add_36383_comb;
  wire [15:0] p1_add_36384_comb;
  wire [15:0] p1_add_36391_comb;
  wire [15:0] p1_add_36392_comb;
  wire [15:0] p1_add_36393_comb;
  wire [15:0] p1_add_36399_comb;
  wire [15:0] p1_add_36400_comb;
  wire [15:0] p1_add_36401_comb;
  wire [15:0] p1_add_36402_comb;
  wire [15:0] p1_add_36407_comb;
  wire [15:0] p1_add_36408_comb;
  wire [15:0] p1_add_36409_comb;
  wire [15:0] p1_add_36410_comb;
  wire [15:0] p1_add_36411_comb;
  wire [15:0] p1_add_36415_comb;
  wire [15:0] p1_add_36416_comb;
  wire [15:0] p1_add_36417_comb;
  wire [15:0] p1_add_36418_comb;
  wire [15:0] p1_add_36419_comb;
  wire [15:0] p1_add_36420_comb;
  wire [15:0] p1_add_36423_comb;
  wire [15:0] p1_add_36424_comb;
  wire [15:0] p1_add_36425_comb;
  wire [15:0] p1_add_36426_comb;
  wire [15:0] p1_add_36427_comb;
  wire [15:0] p1_add_36428_comb;
  wire [15:0] p1_add_36429_comb;
  wire [15:0] p1_add_36431_comb;
  wire [15:0] p1_add_36432_comb;
  wire [15:0] p1_add_36433_comb;
  wire [15:0] p1_add_36434_comb;
  wire [15:0] p1_add_36435_comb;
  wire [15:0] p1_add_36436_comb;
  wire [15:0] p1_add_36437_comb;
  wire [15:0] p1_add_36438_comb;
  wire [31:0] p1_smul_36439_comb;
  wire [31:0] p1_smul_36440_comb;
  wire [31:0] p1_smul_36443_comb;
  wire [15:0] p1_add_36448_comb;
  wire [15:0] p1_add_36452_comb;
  wire [15:0] p1_add_36453_comb;
  wire [15:0] p1_add_36456_comb;
  wire [15:0] p1_add_36457_comb;
  wire [15:0] p1_add_36458_comb;
  wire [15:0] p1_add_36460_comb;
  wire [15:0] p1_add_36461_comb;
  wire [15:0] p1_add_36462_comb;
  wire [15:0] p1_add_36463_comb;
  wire [15:0] p1_add_36464_comb;
  wire [15:0] p1_add_36465_comb;
  wire [15:0] p1_add_36466_comb;
  wire [15:0] p1_add_36467_comb;
  wire [15:0] p1_add_36468_comb;
  wire [15:0] p1_add_36469_comb;
  wire [15:0] p1_add_36470_comb;
  wire [15:0] p1_add_36471_comb;
  wire [15:0] p1_add_36472_comb;
  wire [15:0] p1_add_36473_comb;
  wire [15:0] p1_add_36474_comb;
  wire [15:0] p1_add_36475_comb;
  wire [15:0] p1_add_36476_comb;
  wire [15:0] p1_add_36477_comb;
  wire [15:0] p1_add_36478_comb;
  wire [15:0] p1_add_36479_comb;
  wire [15:0] p1_add_36480_comb;
  wire [15:0] p1_add_36481_comb;
  wire [15:0] p1_add_36482_comb;
  wire [15:0] p1_add_36483_comb;
  wire [15:0] p1_add_36484_comb;
  wire [15:0] p1_add_36485_comb;
  wire [15:0] p1_add_36486_comb;
  wire [15:0] p1_add_36487_comb;
  wire [15:0] p1_add_36488_comb;
  wire [15:0] p1_add_36489_comb;
  wire [15:0] p1_add_36490_comb;
  wire [15:0] p1_add_36491_comb;
  wire [15:0] p1_add_36492_comb;
  wire [15:0] p1_add_36493_comb;
  wire [15:0] p1_add_36494_comb;
  wire [15:0] p1_add_36495_comb;
  wire [31:0] p1_smul_36496_comb;
  wire [15:0] p1_add_36499_comb;
  wire [15:0] p1_add_36501_comb;
  wire [15:0] p1_add_36502_comb;
  wire [15:0] p1_add_36503_comb;
  wire [15:0] p1_add_36504_comb;
  wire [15:0] p1_add_36505_comb;
  wire [15:0] p1_add_36506_comb;
  wire [15:0] p1_add_36507_comb;
  wire [15:0] p1_add_36508_comb;
  wire [15:0] p1_add_36509_comb;
  wire [15:0] p1_add_36510_comb;
  wire [15:0] p1_add_36511_comb;
  wire [15:0] p1_add_36512_comb;
  wire [15:0] p1_add_36513_comb;
  wire [15:0] p1_add_36514_comb;
  wire [15:0] p1_add_36515_comb;
  wire [15:0] p1_add_36516_comb;
  wire [15:0] p1_add_36517_comb;
  wire [15:0] p1_add_36518_comb;
  wire [15:0] p1_add_36519_comb;
  wire [15:0] p1_add_36520_comb;
  wire [15:0] p1_add_36521_comb;
  wire [15:0] p1_add_36522_comb;
  wire [15:0] p1_add_36523_comb;
  wire [15:0] p1_add_36524_comb;
  wire [15:0] p1_add_36525_comb;
  wire [15:0] p1_add_36526_comb;
  wire [15:0] p1_add_36528_comb;
  wire [15:0] p1_add_36529_comb;
  wire [15:0] p1_add_36530_comb;
  wire [15:0] p1_add_36531_comb;
  wire [15:0] p1_add_36532_comb;
  wire [15:0] p1_add_36533_comb;
  wire [15:0] p1_add_36534_comb;
  wire [15:0] p1_add_36535_comb;
  wire [15:0] p1_add_36536_comb;
  wire [15:0] p1_add_36537_comb;
  wire [15:0] p1_add_36538_comb;
  wire [15:0] p1_add_36539_comb;
  wire [15:0] p1_add_36540_comb;
  wire [15:0] p1_add_36541_comb;
  wire [15:0] p1_add_36542_comb;
  wire [15:0] p1_neg_36543_comb;
  wire [15:0] p1_neg_36544_comb;
  wire [15:0] p1_neg_36545_comb;
  wire [15:0] p1_neg_36546_comb;
  wire [15:0] p1_neg_36547_comb;
  wire [15:0] p1_neg_36548_comb;
  wire [15:0] p1_neg_36549_comb;
  wire [15:0] p1_neg_36550_comb;
  wire [15:0] p1_neg_36551_comb;
  wire [15:0] p1_neg_36552_comb;
  wire [15:0] p1_neg_36553_comb;
  wire [15:0] p1_neg_36554_comb;
  wire [15:0] p1_neg_36555_comb;
  wire [15:0] p1_neg_36556_comb;
  wire [15:0] p1_neg_36557_comb;
  wire [15:0] p1_neg_36558_comb;
  wire [31:0] p1_sign_ext_36559_comb;
  wire [31:0] p1_sign_ext_36560_comb;
  wire [31:0] p1_sign_ext_36561_comb;
  wire [31:0] p1_sign_ext_36562_comb;
  wire [31:0] p1_sign_ext_36563_comb;
  wire [31:0] p1_sign_ext_36564_comb;
  wire [31:0] p1_sign_ext_36565_comb;
  wire [31:0] p1_sign_ext_36566_comb;
  assign p1_array_index_36119_comb = p0_signal[4'h8];
  assign p1_array_index_36120_comb = p0_kernel[4'h0];
  assign p1_array_index_36121_comb = p0_signal[4'h7];
  assign p1_array_index_36122_comb = p0_kernel[4'h1];
  assign p1_array_index_36123_comb = p0_signal[4'h9];
  assign p1_array_index_36124_comb = p0_kernel[4'h2];
  assign p1_array_index_36125_comb = p0_signal[4'h6];
  assign p1_array_index_36126_comb = p0_kernel[4'h3];
  assign p1_array_index_36127_comb = p0_signal[4'ha];
  assign p1_array_index_36128_comb = p0_kernel[4'h4];
  assign p1_array_index_36129_comb = p0_signal[4'h5];
  assign p1_array_index_36130_comb = p0_kernel[4'h5];
  assign p1_array_index_36131_comb = p0_signal[4'hb];
  assign p1_array_index_36132_comb = p0_kernel[4'h6];
  assign p1_array_index_36133_comb = p0_signal[4'h4];
  assign p1_array_index_36134_comb = p0_kernel[4'h7];
  assign p1_array_index_36135_comb = p0_signal[4'hc];
  assign p1_array_index_36136_comb = p0_kernel[4'h8];
  assign p1_array_index_36137_comb = p0_signal[4'h3];
  assign p1_array_index_36138_comb = p0_kernel[4'h9];
  assign p1_array_index_36139_comb = p0_signal[4'hd];
  assign p1_array_index_36140_comb = p0_kernel[4'ha];
  assign p1_array_index_36141_comb = p0_signal[4'h2];
  assign p1_array_index_36142_comb = p0_kernel[4'hb];
  assign p1_array_index_36143_comb = p0_signal[4'he];
  assign p1_array_index_36144_comb = p0_kernel[4'hc];
  assign p1_array_index_36145_comb = p0_signal[4'h1];
  assign p1_array_index_36146_comb = p0_kernel[4'hd];
  assign p1_array_index_36148_comb = p0_kernel[4'he];
  assign p1_array_index_36149_comb = p0_signal[4'h0];
  assign p1_smul_36151_comb = smul32b_16b_x_16b(p1_array_index_36119_comb, p1_array_index_36120_comb);
  assign p1_smul_36152_comb = smul32b_16b_x_16b(p1_array_index_36121_comb, p1_array_index_36122_comb);
  assign p1_smul_36153_comb = smul32b_16b_x_16b(p1_array_index_36123_comb, p1_array_index_36120_comb);
  assign p1_smul_36154_comb = smul32b_16b_x_16b(p1_array_index_36119_comb, p1_array_index_36122_comb);
  assign p1_smul_36155_comb = smul32b_16b_x_16b(p1_array_index_36121_comb, p1_array_index_36124_comb);
  assign p1_smul_36156_comb = smul32b_16b_x_16b(p1_array_index_36125_comb, p1_array_index_36126_comb);
  assign p1_smul_36157_comb = smul32b_16b_x_16b(p1_array_index_36127_comb, p1_array_index_36120_comb);
  assign p1_smul_36158_comb = smul32b_16b_x_16b(p1_array_index_36123_comb, p1_array_index_36122_comb);
  assign p1_smul_36159_comb = smul32b_16b_x_16b(p1_array_index_36119_comb, p1_array_index_36124_comb);
  assign p1_smul_36160_comb = smul32b_16b_x_16b(p1_array_index_36121_comb, p1_array_index_36126_comb);
  assign p1_smul_36161_comb = smul32b_16b_x_16b(p1_array_index_36125_comb, p1_array_index_36128_comb);
  assign p1_smul_36162_comb = smul32b_16b_x_16b(p1_array_index_36129_comb, p1_array_index_36130_comb);
  assign p1_smul_36163_comb = smul32b_16b_x_16b(p1_array_index_36131_comb, p1_array_index_36120_comb);
  assign p1_smul_36164_comb = smul32b_16b_x_16b(p1_array_index_36127_comb, p1_array_index_36122_comb);
  assign p1_smul_36165_comb = smul32b_16b_x_16b(p1_array_index_36123_comb, p1_array_index_36124_comb);
  assign p1_smul_36166_comb = smul32b_16b_x_16b(p1_array_index_36119_comb, p1_array_index_36126_comb);
  assign p1_smul_36167_comb = smul32b_16b_x_16b(p1_array_index_36121_comb, p1_array_index_36128_comb);
  assign p1_smul_36168_comb = smul32b_16b_x_16b(p1_array_index_36125_comb, p1_array_index_36130_comb);
  assign p1_smul_36169_comb = smul32b_16b_x_16b(p1_array_index_36129_comb, p1_array_index_36132_comb);
  assign p1_smul_36170_comb = smul32b_16b_x_16b(p1_array_index_36133_comb, p1_array_index_36134_comb);
  assign p1_smul_36171_comb = smul32b_16b_x_16b(p1_array_index_36135_comb, p1_array_index_36120_comb);
  assign p1_smul_36172_comb = smul32b_16b_x_16b(p1_array_index_36131_comb, p1_array_index_36122_comb);
  assign p1_smul_36173_comb = smul32b_16b_x_16b(p1_array_index_36127_comb, p1_array_index_36124_comb);
  assign p1_smul_36174_comb = smul32b_16b_x_16b(p1_array_index_36123_comb, p1_array_index_36126_comb);
  assign p1_smul_36175_comb = smul32b_16b_x_16b(p1_array_index_36119_comb, p1_array_index_36128_comb);
  assign p1_smul_36176_comb = smul32b_16b_x_16b(p1_array_index_36121_comb, p1_array_index_36130_comb);
  assign p1_smul_36177_comb = smul32b_16b_x_16b(p1_array_index_36125_comb, p1_array_index_36132_comb);
  assign p1_smul_36178_comb = smul32b_16b_x_16b(p1_array_index_36129_comb, p1_array_index_36134_comb);
  assign p1_smul_36179_comb = smul32b_16b_x_16b(p1_array_index_36133_comb, p1_array_index_36136_comb);
  assign p1_smul_36180_comb = smul32b_16b_x_16b(p1_array_index_36137_comb, p1_array_index_36138_comb);
  assign p1_smul_36181_comb = smul32b_16b_x_16b(p1_array_index_36139_comb, p1_array_index_36120_comb);
  assign p1_smul_36182_comb = smul32b_16b_x_16b(p1_array_index_36135_comb, p1_array_index_36122_comb);
  assign p1_smul_36183_comb = smul32b_16b_x_16b(p1_array_index_36131_comb, p1_array_index_36124_comb);
  assign p1_smul_36184_comb = smul32b_16b_x_16b(p1_array_index_36127_comb, p1_array_index_36126_comb);
  assign p1_smul_36185_comb = smul32b_16b_x_16b(p1_array_index_36123_comb, p1_array_index_36128_comb);
  assign p1_smul_36186_comb = smul32b_16b_x_16b(p1_array_index_36119_comb, p1_array_index_36130_comb);
  assign p1_smul_36187_comb = smul32b_16b_x_16b(p1_array_index_36121_comb, p1_array_index_36132_comb);
  assign p1_smul_36188_comb = smul32b_16b_x_16b(p1_array_index_36125_comb, p1_array_index_36134_comb);
  assign p1_smul_36189_comb = smul32b_16b_x_16b(p1_array_index_36129_comb, p1_array_index_36136_comb);
  assign p1_smul_36190_comb = smul32b_16b_x_16b(p1_array_index_36133_comb, p1_array_index_36138_comb);
  assign p1_smul_36191_comb = smul32b_16b_x_16b(p1_array_index_36137_comb, p1_array_index_36140_comb);
  assign p1_smul_36192_comb = smul32b_16b_x_16b(p1_array_index_36141_comb, p1_array_index_36142_comb);
  assign p1_smul_36193_comb = smul32b_16b_x_16b(p1_array_index_36143_comb, p1_array_index_36120_comb);
  assign p1_smul_36194_comb = smul32b_16b_x_16b(p1_array_index_36139_comb, p1_array_index_36122_comb);
  assign p1_smul_36195_comb = smul32b_16b_x_16b(p1_array_index_36135_comb, p1_array_index_36124_comb);
  assign p1_smul_36196_comb = smul32b_16b_x_16b(p1_array_index_36131_comb, p1_array_index_36126_comb);
  assign p1_smul_36197_comb = smul32b_16b_x_16b(p1_array_index_36127_comb, p1_array_index_36128_comb);
  assign p1_smul_36198_comb = smul32b_16b_x_16b(p1_array_index_36123_comb, p1_array_index_36130_comb);
  assign p1_smul_36199_comb = smul32b_16b_x_16b(p1_array_index_36119_comb, p1_array_index_36132_comb);
  assign p1_smul_36200_comb = smul32b_16b_x_16b(p1_array_index_36121_comb, p1_array_index_36134_comb);
  assign p1_smul_36201_comb = smul32b_16b_x_16b(p1_array_index_36125_comb, p1_array_index_36136_comb);
  assign p1_smul_36202_comb = smul32b_16b_x_16b(p1_array_index_36129_comb, p1_array_index_36138_comb);
  assign p1_smul_36203_comb = smul32b_16b_x_16b(p1_array_index_36133_comb, p1_array_index_36140_comb);
  assign p1_smul_36204_comb = smul32b_16b_x_16b(p1_array_index_36137_comb, p1_array_index_36142_comb);
  assign p1_smul_36205_comb = smul32b_16b_x_16b(p1_array_index_36141_comb, p1_array_index_36144_comb);
  assign p1_smul_36206_comb = smul32b_16b_x_16b(p1_array_index_36145_comb, p1_array_index_36146_comb);
  assign p1_smul_36207_comb = smul32b_16b_x_16b(p0_signal[4'hf], p1_array_index_36120_comb);
  assign p1_smul_36208_comb = smul32b_16b_x_16b(p1_array_index_36143_comb, p1_array_index_36122_comb);
  assign p1_smul_36209_comb = smul32b_16b_x_16b(p1_array_index_36139_comb, p1_array_index_36124_comb);
  assign p1_smul_36210_comb = smul32b_16b_x_16b(p1_array_index_36135_comb, p1_array_index_36126_comb);
  assign p1_smul_36211_comb = smul32b_16b_x_16b(p1_array_index_36131_comb, p1_array_index_36128_comb);
  assign p1_smul_36212_comb = smul32b_16b_x_16b(p1_array_index_36127_comb, p1_array_index_36130_comb);
  assign p1_smul_36213_comb = smul32b_16b_x_16b(p1_array_index_36123_comb, p1_array_index_36132_comb);
  assign p1_smul_36214_comb = smul32b_16b_x_16b(p1_array_index_36119_comb, p1_array_index_36134_comb);
  assign p1_smul_36215_comb = smul32b_16b_x_16b(p1_array_index_36121_comb, p1_array_index_36136_comb);
  assign p1_smul_36216_comb = smul32b_16b_x_16b(p1_array_index_36125_comb, p1_array_index_36138_comb);
  assign p1_smul_36217_comb = smul32b_16b_x_16b(p1_array_index_36129_comb, p1_array_index_36140_comb);
  assign p1_smul_36218_comb = smul32b_16b_x_16b(p1_array_index_36133_comb, p1_array_index_36142_comb);
  assign p1_smul_36219_comb = smul32b_16b_x_16b(p1_array_index_36137_comb, p1_array_index_36144_comb);
  assign p1_smul_36220_comb = smul32b_16b_x_16b(p1_array_index_36141_comb, p1_array_index_36146_comb);
  assign p1_smul_36221_comb = smul32b_16b_x_16b(p1_array_index_36145_comb, p1_array_index_36148_comb);
  assign p1_smul_36222_comb = smul32b_16b_x_16b(p1_array_index_36149_comb, p0_kernel[4'hf]);
  assign p1_smul_36223_comb = smul32b_16b_x_16b(p1_array_index_36133_comb, p1_array_index_36120_comb);
  assign p1_smul_36224_comb = smul32b_16b_x_16b(p1_array_index_36137_comb, p1_array_index_36122_comb);
  assign p1_smul_36225_comb = smul32b_16b_x_16b(p1_array_index_36129_comb, p1_array_index_36120_comb);
  assign p1_smul_36226_comb = smul32b_16b_x_16b(p1_array_index_36133_comb, p1_array_index_36122_comb);
  assign p1_smul_36227_comb = smul32b_16b_x_16b(p1_array_index_36137_comb, p1_array_index_36124_comb);
  assign p1_smul_36228_comb = smul32b_16b_x_16b(p1_array_index_36141_comb, p1_array_index_36126_comb);
  assign p1_smul_36229_comb = smul32b_16b_x_16b(p1_array_index_36125_comb, p1_array_index_36120_comb);
  assign p1_smul_36230_comb = smul32b_16b_x_16b(p1_array_index_36129_comb, p1_array_index_36122_comb);
  assign p1_smul_36231_comb = smul32b_16b_x_16b(p1_array_index_36133_comb, p1_array_index_36124_comb);
  assign p1_smul_36232_comb = smul32b_16b_x_16b(p1_array_index_36137_comb, p1_array_index_36126_comb);
  assign p1_smul_36233_comb = smul32b_16b_x_16b(p1_array_index_36141_comb, p1_array_index_36128_comb);
  assign p1_smul_36234_comb = smul32b_16b_x_16b(p1_array_index_36145_comb, p1_array_index_36130_comb);
  assign p1_smul_36235_comb = smul32b_16b_x_16b(p1_array_index_36121_comb, p1_array_index_36120_comb);
  assign p1_smul_36236_comb = smul32b_16b_x_16b(p1_array_index_36125_comb, p1_array_index_36122_comb);
  assign p1_smul_36237_comb = smul32b_16b_x_16b(p1_array_index_36129_comb, p1_array_index_36124_comb);
  assign p1_smul_36238_comb = smul32b_16b_x_16b(p1_array_index_36133_comb, p1_array_index_36126_comb);
  assign p1_smul_36239_comb = smul32b_16b_x_16b(p1_array_index_36137_comb, p1_array_index_36128_comb);
  assign p1_smul_36240_comb = smul32b_16b_x_16b(p1_array_index_36141_comb, p1_array_index_36130_comb);
  assign p1_smul_36241_comb = smul32b_16b_x_16b(p1_array_index_36145_comb, p1_array_index_36132_comb);
  assign p1_smul_36242_comb = smul32b_16b_x_16b(p1_array_index_36149_comb, p1_array_index_36134_comb);
  assign p1_smul_36245_comb = smul32b_16b_x_16b(p1_array_index_36125_comb, p1_array_index_36124_comb);
  assign p1_smul_36246_comb = smul32b_16b_x_16b(p1_array_index_36129_comb, p1_array_index_36126_comb);
  assign p1_smul_36247_comb = smul32b_16b_x_16b(p1_array_index_36133_comb, p1_array_index_36128_comb);
  assign p1_smul_36248_comb = smul32b_16b_x_16b(p1_array_index_36137_comb, p1_array_index_36130_comb);
  assign p1_smul_36249_comb = smul32b_16b_x_16b(p1_array_index_36141_comb, p1_array_index_36132_comb);
  assign p1_smul_36250_comb = smul32b_16b_x_16b(p1_array_index_36145_comb, p1_array_index_36134_comb);
  assign p1_smul_36251_comb = smul32b_16b_x_16b(p1_array_index_36149_comb, p1_array_index_36136_comb);
  assign p1_smul_36256_comb = smul32b_16b_x_16b(p1_array_index_36129_comb, p1_array_index_36128_comb);
  assign p1_smul_36257_comb = smul32b_16b_x_16b(p1_array_index_36133_comb, p1_array_index_36130_comb);
  assign p1_smul_36258_comb = smul32b_16b_x_16b(p1_array_index_36137_comb, p1_array_index_36132_comb);
  assign p1_smul_36259_comb = smul32b_16b_x_16b(p1_array_index_36141_comb, p1_array_index_36134_comb);
  assign p1_smul_36260_comb = smul32b_16b_x_16b(p1_array_index_36145_comb, p1_array_index_36136_comb);
  assign p1_smul_36261_comb = smul32b_16b_x_16b(p1_array_index_36149_comb, p1_array_index_36138_comb);
  assign p1_smul_36268_comb = smul32b_16b_x_16b(p1_array_index_36133_comb, p1_array_index_36132_comb);
  assign p1_smul_36269_comb = smul32b_16b_x_16b(p1_array_index_36137_comb, p1_array_index_36134_comb);
  assign p1_smul_36270_comb = smul32b_16b_x_16b(p1_array_index_36141_comb, p1_array_index_36136_comb);
  assign p1_smul_36271_comb = smul32b_16b_x_16b(p1_array_index_36145_comb, p1_array_index_36138_comb);
  assign p1_smul_36272_comb = smul32b_16b_x_16b(p1_array_index_36149_comb, p1_array_index_36140_comb);
  assign p1_smul_36281_comb = smul32b_16b_x_16b(p1_array_index_36137_comb, p1_array_index_36136_comb);
  assign p1_smul_36282_comb = smul32b_16b_x_16b(p1_array_index_36141_comb, p1_array_index_36138_comb);
  assign p1_smul_36283_comb = smul32b_16b_x_16b(p1_array_index_36145_comb, p1_array_index_36140_comb);
  assign p1_smul_36284_comb = smul32b_16b_x_16b(p1_array_index_36149_comb, p1_array_index_36142_comb);
  assign p1_smul_36295_comb = smul32b_16b_x_16b(p1_array_index_36141_comb, p1_array_index_36140_comb);
  assign p1_smul_36296_comb = smul32b_16b_x_16b(p1_array_index_36145_comb, p1_array_index_36142_comb);
  assign p1_smul_36297_comb = smul32b_16b_x_16b(p1_array_index_36149_comb, p1_array_index_36144_comb);
  assign p1_smul_36310_comb = smul32b_16b_x_16b(p1_array_index_36145_comb, p1_array_index_36144_comb);
  assign p1_smul_36311_comb = smul32b_16b_x_16b(p1_array_index_36149_comb, p1_array_index_36146_comb);
  assign p1_smul_36326_comb = smul32b_16b_x_16b(p1_array_index_36149_comb, p1_array_index_36148_comb);
  assign p1_smul_36343_comb = smul32b_16b_x_16b(p1_array_index_36141_comb, p1_array_index_36120_comb);
  assign p1_smul_36344_comb = smul32b_16b_x_16b(p1_array_index_36145_comb, p1_array_index_36122_comb);
  assign p1_smul_36345_comb = smul32b_16b_x_16b(p1_array_index_36137_comb, p1_array_index_36120_comb);
  assign p1_smul_36346_comb = smul32b_16b_x_16b(p1_array_index_36141_comb, p1_array_index_36122_comb);
  assign p1_smul_36347_comb = smul32b_16b_x_16b(p1_array_index_36145_comb, p1_array_index_36124_comb);
  assign p1_smul_36348_comb = smul32b_16b_x_16b(p1_array_index_36149_comb, p1_array_index_36126_comb);
  assign p1_smul_36351_comb = smul32b_16b_x_16b(p1_array_index_36141_comb, p1_array_index_36124_comb);
  assign p1_smul_36352_comb = smul32b_16b_x_16b(p1_array_index_36145_comb, p1_array_index_36126_comb);
  assign p1_smul_36353_comb = smul32b_16b_x_16b(p1_array_index_36149_comb, p1_array_index_36128_comb);
  assign p1_smul_36358_comb = smul32b_16b_x_16b(p1_array_index_36145_comb, p1_array_index_36128_comb);
  assign p1_smul_36359_comb = smul32b_16b_x_16b(p1_array_index_36149_comb, p1_array_index_36130_comb);
  assign p1_smul_36366_comb = smul32b_16b_x_16b(p1_array_index_36149_comb, p1_array_index_36132_comb);
  assign p1_add_36375_comb = p1_smul_36151_comb[15:0] + p1_smul_36152_comb[15:0];
  assign p1_add_36383_comb = p1_smul_36153_comb[15:0] + p1_smul_36154_comb[15:0];
  assign p1_add_36384_comb = p1_smul_36155_comb[15:0] + p1_smul_36156_comb[15:0];
  assign p1_add_36391_comb = p1_smul_36157_comb[15:0] + p1_smul_36158_comb[15:0];
  assign p1_add_36392_comb = p1_smul_36159_comb[15:0] + p1_smul_36160_comb[15:0];
  assign p1_add_36393_comb = p1_smul_36161_comb[15:0] + p1_smul_36162_comb[15:0];
  assign p1_add_36399_comb = p1_smul_36163_comb[15:0] + p1_smul_36164_comb[15:0];
  assign p1_add_36400_comb = p1_smul_36165_comb[15:0] + p1_smul_36166_comb[15:0];
  assign p1_add_36401_comb = p1_smul_36167_comb[15:0] + p1_smul_36168_comb[15:0];
  assign p1_add_36402_comb = p1_smul_36169_comb[15:0] + p1_smul_36170_comb[15:0];
  assign p1_add_36407_comb = p1_smul_36171_comb[15:0] + p1_smul_36172_comb[15:0];
  assign p1_add_36408_comb = p1_smul_36173_comb[15:0] + p1_smul_36174_comb[15:0];
  assign p1_add_36409_comb = p1_smul_36175_comb[15:0] + p1_smul_36176_comb[15:0];
  assign p1_add_36410_comb = p1_smul_36177_comb[15:0] + p1_smul_36178_comb[15:0];
  assign p1_add_36411_comb = p1_smul_36179_comb[15:0] + p1_smul_36180_comb[15:0];
  assign p1_add_36415_comb = p1_smul_36181_comb[15:0] + p1_smul_36182_comb[15:0];
  assign p1_add_36416_comb = p1_smul_36183_comb[15:0] + p1_smul_36184_comb[15:0];
  assign p1_add_36417_comb = p1_smul_36185_comb[15:0] + p1_smul_36186_comb[15:0];
  assign p1_add_36418_comb = p1_smul_36187_comb[15:0] + p1_smul_36188_comb[15:0];
  assign p1_add_36419_comb = p1_smul_36189_comb[15:0] + p1_smul_36190_comb[15:0];
  assign p1_add_36420_comb = p1_smul_36191_comb[15:0] + p1_smul_36192_comb[15:0];
  assign p1_add_36423_comb = p1_smul_36193_comb[15:0] + p1_smul_36194_comb[15:0];
  assign p1_add_36424_comb = p1_smul_36195_comb[15:0] + p1_smul_36196_comb[15:0];
  assign p1_add_36425_comb = p1_smul_36197_comb[15:0] + p1_smul_36198_comb[15:0];
  assign p1_add_36426_comb = p1_smul_36199_comb[15:0] + p1_smul_36200_comb[15:0];
  assign p1_add_36427_comb = p1_smul_36201_comb[15:0] + p1_smul_36202_comb[15:0];
  assign p1_add_36428_comb = p1_smul_36203_comb[15:0] + p1_smul_36204_comb[15:0];
  assign p1_add_36429_comb = p1_smul_36205_comb[15:0] + p1_smul_36206_comb[15:0];
  assign p1_add_36431_comb = p1_smul_36207_comb[15:0] + p1_smul_36208_comb[15:0];
  assign p1_add_36432_comb = p1_smul_36209_comb[15:0] + p1_smul_36210_comb[15:0];
  assign p1_add_36433_comb = p1_smul_36211_comb[15:0] + p1_smul_36212_comb[15:0];
  assign p1_add_36434_comb = p1_smul_36213_comb[15:0] + p1_smul_36214_comb[15:0];
  assign p1_add_36435_comb = p1_smul_36215_comb[15:0] + p1_smul_36216_comb[15:0];
  assign p1_add_36436_comb = p1_smul_36217_comb[15:0] + p1_smul_36218_comb[15:0];
  assign p1_add_36437_comb = p1_smul_36219_comb[15:0] + p1_smul_36220_comb[15:0];
  assign p1_add_36438_comb = p1_smul_36221_comb[15:0] + p1_smul_36222_comb[15:0];
  assign p1_smul_36439_comb = smul32b_16b_x_16b(p1_array_index_36145_comb, p1_array_index_36120_comb);
  assign p1_smul_36440_comb = smul32b_16b_x_16b(p1_array_index_36149_comb, p1_array_index_36122_comb);
  assign p1_smul_36443_comb = smul32b_16b_x_16b(p1_array_index_36149_comb, p1_array_index_36124_comb);
  assign p1_add_36448_comb = p1_smul_36223_comb[15:0] + p1_smul_36224_comb[15:0];
  assign p1_add_36452_comb = p1_smul_36225_comb[15:0] + p1_smul_36226_comb[15:0];
  assign p1_add_36453_comb = p1_smul_36227_comb[15:0] + p1_smul_36228_comb[15:0];
  assign p1_add_36456_comb = p1_smul_36229_comb[15:0] + p1_smul_36230_comb[15:0];
  assign p1_add_36457_comb = p1_smul_36231_comb[15:0] + p1_smul_36232_comb[15:0];
  assign p1_add_36458_comb = p1_smul_36233_comb[15:0] + p1_smul_36234_comb[15:0];
  assign p1_add_36460_comb = p1_smul_36235_comb[15:0] + p1_smul_36236_comb[15:0];
  assign p1_add_36461_comb = p1_smul_36237_comb[15:0] + p1_smul_36238_comb[15:0];
  assign p1_add_36462_comb = p1_smul_36239_comb[15:0] + p1_smul_36240_comb[15:0];
  assign p1_add_36463_comb = p1_smul_36241_comb[15:0] + p1_smul_36242_comb[15:0];
  assign p1_add_36464_comb = p1_add_36375_comb + p1_smul_36245_comb[15:0];
  assign p1_add_36465_comb = p1_smul_36246_comb[15:0] + p1_smul_36247_comb[15:0];
  assign p1_add_36466_comb = p1_smul_36248_comb[15:0] + p1_smul_36249_comb[15:0];
  assign p1_add_36467_comb = p1_smul_36250_comb[15:0] + p1_smul_36251_comb[15:0];
  assign p1_add_36468_comb = p1_add_36383_comb + p1_add_36384_comb;
  assign p1_add_36469_comb = p1_smul_36256_comb[15:0] + p1_smul_36257_comb[15:0];
  assign p1_add_36470_comb = p1_smul_36258_comb[15:0] + p1_smul_36259_comb[15:0];
  assign p1_add_36471_comb = p1_smul_36260_comb[15:0] + p1_smul_36261_comb[15:0];
  assign p1_add_36472_comb = p1_add_36391_comb + p1_add_36392_comb;
  assign p1_add_36473_comb = p1_add_36393_comb + p1_smul_36268_comb[15:0];
  assign p1_add_36474_comb = p1_smul_36269_comb[15:0] + p1_smul_36270_comb[15:0];
  assign p1_add_36475_comb = p1_smul_36271_comb[15:0] + p1_smul_36272_comb[15:0];
  assign p1_add_36476_comb = p1_add_36399_comb + p1_add_36400_comb;
  assign p1_add_36477_comb = p1_add_36401_comb + p1_add_36402_comb;
  assign p1_add_36478_comb = p1_smul_36281_comb[15:0] + p1_smul_36282_comb[15:0];
  assign p1_add_36479_comb = p1_smul_36283_comb[15:0] + p1_smul_36284_comb[15:0];
  assign p1_add_36480_comb = p1_add_36407_comb + p1_add_36408_comb;
  assign p1_add_36481_comb = p1_add_36409_comb + p1_add_36410_comb;
  assign p1_add_36482_comb = p1_add_36411_comb + p1_smul_36295_comb[15:0];
  assign p1_add_36483_comb = p1_smul_36296_comb[15:0] + p1_smul_36297_comb[15:0];
  assign p1_add_36484_comb = p1_add_36415_comb + p1_add_36416_comb;
  assign p1_add_36485_comb = p1_add_36417_comb + p1_add_36418_comb;
  assign p1_add_36486_comb = p1_add_36419_comb + p1_add_36420_comb;
  assign p1_add_36487_comb = p1_smul_36310_comb[15:0] + p1_smul_36311_comb[15:0];
  assign p1_add_36488_comb = p1_add_36423_comb + p1_add_36424_comb;
  assign p1_add_36489_comb = p1_add_36425_comb + p1_add_36426_comb;
  assign p1_add_36490_comb = p1_add_36427_comb + p1_add_36428_comb;
  assign p1_add_36491_comb = p1_add_36429_comb + p1_smul_36326_comb[15:0];
  assign p1_add_36492_comb = p1_add_36431_comb + p1_add_36432_comb;
  assign p1_add_36493_comb = p1_add_36433_comb + p1_add_36434_comb;
  assign p1_add_36494_comb = p1_add_36435_comb + p1_add_36436_comb;
  assign p1_add_36495_comb = p1_add_36437_comb + p1_add_36438_comb;
  assign p1_smul_36496_comb = smul32b_16b_x_16b(p1_array_index_36149_comb, p1_array_index_36120_comb);
  assign p1_add_36499_comb = p1_smul_36343_comb[15:0] + p1_smul_36344_comb[15:0];
  assign p1_add_36501_comb = p1_smul_36345_comb[15:0] + p1_smul_36346_comb[15:0];
  assign p1_add_36502_comb = p1_smul_36347_comb[15:0] + p1_smul_36348_comb[15:0];
  assign p1_add_36503_comb = p1_add_36448_comb + p1_smul_36351_comb[15:0];
  assign p1_add_36504_comb = p1_smul_36352_comb[15:0] + p1_smul_36353_comb[15:0];
  assign p1_add_36505_comb = p1_add_36452_comb + p1_add_36453_comb;
  assign p1_add_36506_comb = p1_smul_36358_comb[15:0] + p1_smul_36359_comb[15:0];
  assign p1_add_36507_comb = p1_add_36456_comb + p1_add_36457_comb;
  assign p1_add_36508_comb = p1_add_36458_comb + p1_smul_36366_comb[15:0];
  assign p1_add_36509_comb = p1_add_36460_comb + p1_add_36461_comb;
  assign p1_add_36510_comb = p1_add_36462_comb + p1_add_36463_comb;
  assign p1_add_36511_comb = p1_add_36464_comb + p1_add_36465_comb;
  assign p1_add_36512_comb = p1_add_36466_comb + p1_add_36467_comb;
  assign p1_add_36513_comb = p1_add_36468_comb + p1_add_36469_comb;
  assign p1_add_36514_comb = p1_add_36470_comb + p1_add_36471_comb;
  assign p1_add_36515_comb = p1_add_36472_comb + p1_add_36473_comb;
  assign p1_add_36516_comb = p1_add_36474_comb + p1_add_36475_comb;
  assign p1_add_36517_comb = p1_add_36476_comb + p1_add_36477_comb;
  assign p1_add_36518_comb = p1_add_36478_comb + p1_add_36479_comb;
  assign p1_add_36519_comb = p1_add_36480_comb + p1_add_36481_comb;
  assign p1_add_36520_comb = p1_add_36482_comb + p1_add_36483_comb;
  assign p1_add_36521_comb = p1_add_36484_comb + p1_add_36485_comb;
  assign p1_add_36522_comb = p1_add_36486_comb + p1_add_36487_comb;
  assign p1_add_36523_comb = p1_add_36488_comb + p1_add_36489_comb;
  assign p1_add_36524_comb = p1_add_36490_comb + p1_add_36491_comb;
  assign p1_add_36525_comb = p1_add_36492_comb + p1_add_36493_comb;
  assign p1_add_36526_comb = p1_add_36494_comb + p1_add_36495_comb;
  assign p1_add_36528_comb = p1_smul_36439_comb[15:0] + p1_smul_36440_comb[15:0];
  assign p1_add_36529_comb = p1_add_36499_comb + p1_smul_36443_comb[15:0];
  assign p1_add_36530_comb = p1_add_36501_comb + p1_add_36502_comb;
  assign p1_add_36531_comb = p1_add_36503_comb + p1_add_36504_comb;
  assign p1_add_36532_comb = p1_add_36505_comb + p1_add_36506_comb;
  assign p1_add_36533_comb = p1_add_36507_comb + p1_add_36508_comb;
  assign p1_add_36534_comb = p1_add_36509_comb + p1_add_36510_comb;
  assign p1_add_36535_comb = p1_add_36511_comb + p1_add_36512_comb;
  assign p1_add_36536_comb = p1_add_36513_comb + p1_add_36514_comb;
  assign p1_add_36537_comb = p1_add_36515_comb + p1_add_36516_comb;
  assign p1_add_36538_comb = p1_add_36517_comb + p1_add_36518_comb;
  assign p1_add_36539_comb = p1_add_36519_comb + p1_add_36520_comb;
  assign p1_add_36540_comb = p1_add_36521_comb + p1_add_36522_comb;
  assign p1_add_36541_comb = p1_add_36523_comb + p1_add_36524_comb;
  assign p1_add_36542_comb = p1_add_36525_comb + p1_add_36526_comb;
  assign p1_neg_36543_comb = -p1_smul_36496_comb[15:0];
  assign p1_neg_36544_comb = -p1_add_36528_comb;
  assign p1_neg_36545_comb = -p1_add_36529_comb;
  assign p1_neg_36546_comb = -p1_add_36530_comb;
  assign p1_neg_36547_comb = -p1_add_36531_comb;
  assign p1_neg_36548_comb = -p1_add_36532_comb;
  assign p1_neg_36549_comb = -p1_add_36533_comb;
  assign p1_neg_36550_comb = -p1_add_36534_comb;
  assign p1_neg_36551_comb = -p1_add_36535_comb;
  assign p1_neg_36552_comb = -p1_add_36536_comb;
  assign p1_neg_36553_comb = -p1_add_36537_comb;
  assign p1_neg_36554_comb = -p1_add_36538_comb;
  assign p1_neg_36555_comb = -p1_add_36539_comb;
  assign p1_neg_36556_comb = -p1_add_36540_comb;
  assign p1_neg_36557_comb = -p1_add_36541_comb;
  assign p1_neg_36558_comb = -p1_add_36542_comb;
  assign p1_sign_ext_36559_comb = {{16{p1_neg_36543_comb[15]}}, p1_neg_36543_comb};
  assign p1_sign_ext_36560_comb = {{16{p1_neg_36544_comb[15]}}, p1_neg_36544_comb};
  assign p1_sign_ext_36561_comb = {{16{p1_neg_36545_comb[15]}}, p1_neg_36545_comb};
  assign p1_sign_ext_36562_comb = {{16{p1_neg_36546_comb[15]}}, p1_neg_36546_comb};
  assign p1_sign_ext_36563_comb = {{16{p1_neg_36547_comb[15]}}, p1_neg_36547_comb};
  assign p1_sign_ext_36564_comb = {{16{p1_neg_36548_comb[15]}}, p1_neg_36548_comb};
  assign p1_sign_ext_36565_comb = {{16{p1_neg_36549_comb[15]}}, p1_neg_36549_comb};
  assign p1_sign_ext_36566_comb = {{16{p1_neg_36550_comb[15]}}, p1_neg_36550_comb};

  // Registers for pipe stage 1:
  reg [15:0] p1_neg_36543;
  reg [15:0] p1_neg_36544;
  reg [15:0] p1_neg_36545;
  reg [15:0] p1_neg_36546;
  reg [15:0] p1_neg_36547;
  reg [15:0] p1_neg_36548;
  reg [15:0] p1_neg_36549;
  reg [15:0] p1_neg_36550;
  reg [15:0] p1_neg_36551;
  reg [15:0] p1_neg_36552;
  reg [15:0] p1_neg_36553;
  reg [15:0] p1_neg_36554;
  reg [15:0] p1_neg_36555;
  reg [15:0] p1_neg_36556;
  reg [15:0] p1_neg_36557;
  reg [15:0] p1_neg_36558;
  reg [31:0] p1_sign_ext_36559;
  reg [31:0] p1_sign_ext_36560;
  reg [31:0] p1_sign_ext_36561;
  reg [31:0] p1_sign_ext_36562;
  reg [31:0] p1_sign_ext_36563;
  reg [31:0] p1_sign_ext_36564;
  reg [31:0] p1_sign_ext_36565;
  reg [31:0] p1_sign_ext_36566;
  always_ff @ (posedge clk) begin
    p1_neg_36543 <= p1_neg_36543_comb;
    p1_neg_36544 <= p1_neg_36544_comb;
    p1_neg_36545 <= p1_neg_36545_comb;
    p1_neg_36546 <= p1_neg_36546_comb;
    p1_neg_36547 <= p1_neg_36547_comb;
    p1_neg_36548 <= p1_neg_36548_comb;
    p1_neg_36549 <= p1_neg_36549_comb;
    p1_neg_36550 <= p1_neg_36550_comb;
    p1_neg_36551 <= p1_neg_36551_comb;
    p1_neg_36552 <= p1_neg_36552_comb;
    p1_neg_36553 <= p1_neg_36553_comb;
    p1_neg_36554 <= p1_neg_36554_comb;
    p1_neg_36555 <= p1_neg_36555_comb;
    p1_neg_36556 <= p1_neg_36556_comb;
    p1_neg_36557 <= p1_neg_36557_comb;
    p1_neg_36558 <= p1_neg_36558_comb;
    p1_sign_ext_36559 <= p1_sign_ext_36559_comb;
    p1_sign_ext_36560 <= p1_sign_ext_36560_comb;
    p1_sign_ext_36561 <= p1_sign_ext_36561_comb;
    p1_sign_ext_36562 <= p1_sign_ext_36562_comb;
    p1_sign_ext_36563 <= p1_sign_ext_36563_comb;
    p1_sign_ext_36564 <= p1_sign_ext_36564_comb;
    p1_sign_ext_36565 <= p1_sign_ext_36565_comb;
    p1_sign_ext_36566 <= p1_sign_ext_36566_comb;
  end

  // ===== Pipe stage 2:
  wire [31:0] p2_sign_ext_36615_comb;
  wire [31:0] p2_sign_ext_36616_comb;
  wire [31:0] p2_sign_ext_36617_comb;
  wire [31:0] p2_sign_ext_36618_comb;
  wire [31:0] p2_sign_ext_36619_comb;
  wire [31:0] p2_sign_ext_36620_comb;
  wire [31:0] p2_sign_ext_36621_comb;
  wire [31:0] p2_sign_ext_36622_comb;
  wire [31:0] p2_add_36687_comb;
  wire [46:0] p2_smul_33601_NarrowedMult__comb;
  wire [31:0] p2_add_36692_comb;
  wire [46:0] p2_smul_33603_NarrowedMult__comb;
  wire [31:0] p2_add_36697_comb;
  wire [46:0] p2_smul_33605_NarrowedMult__comb;
  wire [31:0] p2_add_36702_comb;
  wire [46:0] p2_smul_33607_NarrowedMult__comb;
  wire [31:0] p2_add_36707_comb;
  wire [46:0] p2_smul_33609_NarrowedMult__comb;
  wire [31:0] p2_add_36712_comb;
  wire [46:0] p2_smul_33611_NarrowedMult__comb;
  wire [31:0] p2_add_36717_comb;
  wire [46:0] p2_smul_33613_NarrowedMult__comb;
  wire [31:0] p2_add_36722_comb;
  wire [46:0] p2_smul_33615_NarrowedMult__comb;
  wire [31:0] p2_add_36727_comb;
  wire [46:0] p2_smul_33617_NarrowedMult__comb;
  wire [31:0] p2_add_36732_comb;
  wire [46:0] p2_smul_33619_NarrowedMult__comb;
  wire [31:0] p2_add_36737_comb;
  wire [46:0] p2_smul_33621_NarrowedMult__comb;
  wire [31:0] p2_add_36742_comb;
  wire [46:0] p2_smul_33623_NarrowedMult__comb;
  wire [31:0] p2_add_36747_comb;
  wire [46:0] p2_smul_33625_NarrowedMult__comb;
  wire [31:0] p2_add_36752_comb;
  wire [46:0] p2_smul_33627_NarrowedMult__comb;
  wire [31:0] p2_add_36757_comb;
  wire [46:0] p2_smul_33629_NarrowedMult__comb;
  wire [31:0] p2_add_36762_comb;
  wire [46:0] p2_smul_33631_NarrowedMult__comb;
  wire [15:0] p2_sign_ext_36769_comb;
  wire [47:0] p2_smul_36771_comb;
  wire [15:0] p2_sign_ext_36774_comb;
  wire [47:0] p2_smul_36776_comb;
  wire [15:0] p2_sign_ext_36779_comb;
  wire [47:0] p2_smul_36781_comb;
  wire [15:0] p2_sign_ext_36784_comb;
  wire [47:0] p2_smul_36786_comb;
  wire [15:0] p2_sign_ext_36789_comb;
  wire [47:0] p2_smul_36791_comb;
  wire [15:0] p2_sign_ext_36794_comb;
  wire [47:0] p2_smul_36796_comb;
  wire [15:0] p2_sign_ext_36799_comb;
  wire [47:0] p2_smul_36801_comb;
  wire [15:0] p2_sign_ext_36804_comb;
  wire [47:0] p2_smul_36806_comb;
  wire [15:0] p2_sign_ext_36809_comb;
  wire [47:0] p2_smul_36811_comb;
  wire [15:0] p2_sign_ext_36814_comb;
  wire [47:0] p2_smul_36816_comb;
  wire [15:0] p2_sign_ext_36819_comb;
  wire [47:0] p2_smul_36821_comb;
  wire [15:0] p2_sign_ext_36824_comb;
  wire [47:0] p2_smul_36826_comb;
  wire [15:0] p2_sign_ext_36829_comb;
  wire [47:0] p2_smul_36831_comb;
  wire [15:0] p2_sign_ext_36834_comb;
  wire [47:0] p2_smul_36836_comb;
  wire [15:0] p2_sign_ext_36839_comb;
  wire [47:0] p2_smul_36841_comb;
  wire [15:0] p2_sign_ext_36844_comb;
  wire [47:0] p2_smul_36846_comb;
  wire [15:0] p2_smul_36847_comb;
  wire [15:0] p2_sub_36848_comb;
  wire [31:0] p2_add_36849_comb;
  wire [63:0] p2_sign_ext_36850_comb;
  wire [15:0] p2_smul_36852_comb;
  wire [15:0] p2_sub_36853_comb;
  wire [31:0] p2_add_36854_comb;
  wire [63:0] p2_sign_ext_36855_comb;
  wire [15:0] p2_smul_36857_comb;
  wire [15:0] p2_sub_36858_comb;
  wire [31:0] p2_add_36859_comb;
  wire [63:0] p2_sign_ext_36860_comb;
  wire [15:0] p2_smul_36862_comb;
  wire [15:0] p2_sub_36863_comb;
  wire [31:0] p2_add_36864_comb;
  wire [63:0] p2_sign_ext_36865_comb;
  wire [15:0] p2_smul_36867_comb;
  wire [15:0] p2_sub_36868_comb;
  wire [31:0] p2_add_36869_comb;
  wire [63:0] p2_sign_ext_36870_comb;
  wire [15:0] p2_smul_36872_comb;
  wire [15:0] p2_sub_36873_comb;
  wire [31:0] p2_add_36874_comb;
  wire [63:0] p2_sign_ext_36875_comb;
  wire [15:0] p2_smul_36877_comb;
  wire [15:0] p2_sub_36878_comb;
  wire [31:0] p2_add_36879_comb;
  wire [63:0] p2_sign_ext_36880_comb;
  wire [15:0] p2_smul_36882_comb;
  wire [15:0] p2_sub_36883_comb;
  wire [31:0] p2_add_36884_comb;
  wire [63:0] p2_sign_ext_36885_comb;
  wire [15:0] p2_smul_36887_comb;
  wire [15:0] p2_sub_36888_comb;
  wire [31:0] p2_add_36889_comb;
  wire [63:0] p2_sign_ext_36890_comb;
  wire [15:0] p2_smul_36892_comb;
  wire [15:0] p2_sub_36893_comb;
  wire [31:0] p2_add_36894_comb;
  wire [63:0] p2_sign_ext_36895_comb;
  wire [15:0] p2_smul_36897_comb;
  wire [15:0] p2_sub_36898_comb;
  wire [31:0] p2_add_36899_comb;
  wire [63:0] p2_sign_ext_36900_comb;
  wire [15:0] p2_smul_36902_comb;
  wire [15:0] p2_sub_36903_comb;
  wire [31:0] p2_add_36904_comb;
  wire [63:0] p2_sign_ext_36905_comb;
  wire [15:0] p2_smul_36907_comb;
  wire [15:0] p2_sub_36908_comb;
  wire [31:0] p2_add_36909_comb;
  wire [63:0] p2_sign_ext_36910_comb;
  wire [15:0] p2_smul_36912_comb;
  wire [15:0] p2_sub_36913_comb;
  wire [31:0] p2_add_36914_comb;
  wire [63:0] p2_sign_ext_36915_comb;
  wire [15:0] p2_smul_36917_comb;
  wire [15:0] p2_sub_36918_comb;
  wire [31:0] p2_add_36919_comb;
  wire [63:0] p2_sign_ext_36920_comb;
  wire [15:0] p2_smul_36922_comb;
  wire [15:0] p2_sub_36923_comb;
  wire [31:0] p2_add_36924_comb;
  wire [63:0] p2_sign_ext_36925_comb;
  wire [15:0] p2_smul_36927_comb;
  wire [62:0] p2_sign_ext_36930_comb;
  wire [48:0] p2_smul_36931_comb;
  wire [15:0] p2_smul_36932_comb;
  wire [62:0] p2_sign_ext_36935_comb;
  wire [48:0] p2_smul_36936_comb;
  wire [15:0] p2_smul_36937_comb;
  wire [62:0] p2_sign_ext_36940_comb;
  wire [48:0] p2_smul_36941_comb;
  wire [15:0] p2_smul_36942_comb;
  wire [62:0] p2_sign_ext_36945_comb;
  wire [48:0] p2_smul_36946_comb;
  wire [15:0] p2_smul_36947_comb;
  wire [62:0] p2_sign_ext_36950_comb;
  wire [48:0] p2_smul_36951_comb;
  wire [15:0] p2_smul_36952_comb;
  wire [62:0] p2_sign_ext_36955_comb;
  wire [48:0] p2_smul_36956_comb;
  wire [15:0] p2_smul_36957_comb;
  wire [62:0] p2_sign_ext_36960_comb;
  wire [48:0] p2_smul_36961_comb;
  wire [15:0] p2_smul_36962_comb;
  wire [62:0] p2_sign_ext_36965_comb;
  wire [48:0] p2_smul_36966_comb;
  wire [48:0] p2_smul_36971_comb;
  wire [48:0] p2_smul_36976_comb;
  wire [48:0] p2_smul_36981_comb;
  wire [48:0] p2_smul_36986_comb;
  wire [48:0] p2_smul_36991_comb;
  wire [48:0] p2_smul_36996_comb;
  wire [48:0] p2_smul_37001_comb;
  wire [48:0] p2_smul_37006_comb;
  wire [46:0] p2_smul_37123_comb;
  wire [46:0] p2_smul_37128_comb;
  wire [46:0] p2_smul_37133_comb;
  wire [46:0] p2_smul_37138_comb;
  wire [46:0] p2_smul_37143_comb;
  wire [46:0] p2_smul_37148_comb;
  wire [46:0] p2_smul_37153_comb;
  wire [46:0] p2_smul_37158_comb;
  wire [46:0] p2_smul_37163_comb;
  wire [46:0] p2_smul_37168_comb;
  wire [46:0] p2_smul_37173_comb;
  wire [46:0] p2_smul_37178_comb;
  wire [46:0] p2_smul_37183_comb;
  wire [46:0] p2_smul_37188_comb;
  wire [46:0] p2_smul_37193_comb;
  wire [46:0] p2_smul_37198_comb;
  wire [15:0] p2_smul_36967_comb;
  wire [62:0] p2_sign_ext_36970_comb;
  wire [15:0] p2_smul_36972_comb;
  wire [62:0] p2_sign_ext_36975_comb;
  wire [15:0] p2_smul_36977_comb;
  wire [62:0] p2_sign_ext_36980_comb;
  wire [15:0] p2_smul_36982_comb;
  wire [62:0] p2_sign_ext_36985_comb;
  wire [15:0] p2_smul_36987_comb;
  wire [62:0] p2_sign_ext_36990_comb;
  wire [15:0] p2_smul_36992_comb;
  wire [62:0] p2_sign_ext_36995_comb;
  wire [15:0] p2_smul_36997_comb;
  wire [62:0] p2_sign_ext_37000_comb;
  wire [15:0] p2_smul_37002_comb;
  wire [62:0] p2_sign_ext_37005_comb;
  wire [15:0] p2_smul_37007_comb;
  wire [15:0] p2_sub_37008_comb;
  wire [64:0] p2_sign_ext_37010_comb;
  wire [15:0] p2_smul_37014_comb;
  wire [15:0] p2_sub_37015_comb;
  wire [64:0] p2_sign_ext_37017_comb;
  wire [15:0] p2_smul_37021_comb;
  wire [15:0] p2_sub_37022_comb;
  wire [64:0] p2_sign_ext_37024_comb;
  wire [15:0] p2_smul_37028_comb;
  wire [15:0] p2_sub_37029_comb;
  wire [64:0] p2_sign_ext_37031_comb;
  wire [15:0] p2_smul_37035_comb;
  wire [15:0] p2_sub_37036_comb;
  wire [64:0] p2_sign_ext_37038_comb;
  wire [15:0] p2_smul_37042_comb;
  wire [15:0] p2_sub_37043_comb;
  wire [64:0] p2_sign_ext_37045_comb;
  wire [15:0] p2_smul_37049_comb;
  wire [15:0] p2_sub_37050_comb;
  wire [64:0] p2_sign_ext_37052_comb;
  wire [15:0] p2_smul_37056_comb;
  wire [15:0] p2_sub_37057_comb;
  wire [64:0] p2_sign_ext_37059_comb;
  wire [64:0] p2_sign_ext_37066_comb;
  wire [64:0] p2_sign_ext_37073_comb;
  wire [64:0] p2_sign_ext_37080_comb;
  wire [64:0] p2_sign_ext_37087_comb;
  wire [64:0] p2_sign_ext_37094_comb;
  wire [64:0] p2_sign_ext_37101_comb;
  wire [64:0] p2_sign_ext_37108_comb;
  wire [64:0] p2_sign_ext_37115_comb;
  wire [62:0] p2_sign_ext_37202_comb;
  wire [62:0] p2_sign_ext_37207_comb;
  wire [62:0] p2_sign_ext_37212_comb;
  wire [62:0] p2_sign_ext_37217_comb;
  wire [62:0] p2_sign_ext_37222_comb;
  wire [62:0] p2_sign_ext_37227_comb;
  wire [62:0] p2_sign_ext_37232_comb;
  wire [62:0] p2_sign_ext_37237_comb;
  wire [62:0] p2_sign_ext_37241_comb;
  wire [62:0] p2_sign_ext_37244_comb;
  wire [62:0] p2_sign_ext_37247_comb;
  wire [62:0] p2_sign_ext_37250_comb;
  wire [62:0] p2_sign_ext_37253_comb;
  wire [62:0] p2_sign_ext_37256_comb;
  wire [62:0] p2_sign_ext_37259_comb;
  wire [62:0] p2_sign_ext_37262_comb;
  wire [15:0] p2_smul_37063_comb;
  wire [15:0] p2_sub_37064_comb;
  wire [15:0] p2_smul_37070_comb;
  wire [15:0] p2_sub_37071_comb;
  wire [15:0] p2_smul_37077_comb;
  wire [15:0] p2_sub_37078_comb;
  wire [15:0] p2_smul_37084_comb;
  wire [15:0] p2_sub_37085_comb;
  wire [15:0] p2_smul_37091_comb;
  wire [15:0] p2_sub_37092_comb;
  wire [15:0] p2_smul_37098_comb;
  wire [15:0] p2_sub_37099_comb;
  wire [15:0] p2_smul_37105_comb;
  wire [15:0] p2_sub_37106_comb;
  wire [15:0] p2_smul_37112_comb;
  wire [15:0] p2_sub_37113_comb;
  wire [15:0] p2_smul_37119_comb;
  wire [15:0] p2_sub_37120_comb;
  wire [15:0] p2_smul_37124_comb;
  wire [15:0] p2_sub_37125_comb;
  wire [15:0] p2_smul_37129_comb;
  wire [15:0] p2_sub_37130_comb;
  wire [15:0] p2_smul_37134_comb;
  wire [15:0] p2_sub_37135_comb;
  wire [15:0] p2_smul_37139_comb;
  wire [15:0] p2_sub_37140_comb;
  wire [15:0] p2_smul_37144_comb;
  wire [15:0] p2_sub_37145_comb;
  wire [15:0] p2_smul_37149_comb;
  wire [15:0] p2_sub_37150_comb;
  wire [15:0] p2_smul_37154_comb;
  wire [15:0] p2_sub_37155_comb;
  wire [31:0] p2_add_37201_comb;
  wire [31:0] p2_add_37206_comb;
  wire [31:0] p2_add_37211_comb;
  wire [31:0] p2_add_37216_comb;
  wire [31:0] p2_add_37221_comb;
  wire [31:0] p2_add_37226_comb;
  wire [31:0] p2_add_37231_comb;
  wire [31:0] p2_add_37236_comb;
  wire [31:0] p2_add_37240_comb;
  wire [31:0] p2_add_37243_comb;
  wire [31:0] p2_add_37246_comb;
  wire [31:0] p2_add_37249_comb;
  wire [31:0] p2_add_37252_comb;
  wire [31:0] p2_add_37255_comb;
  wire [31:0] p2_add_37258_comb;
  wire [31:0] p2_add_37261_comb;
  wire [46:0] p2_smul_37265_comb;
  wire [46:0] p2_smul_37268_comb;
  wire [46:0] p2_smul_37271_comb;
  wire [46:0] p2_smul_37274_comb;
  wire [46:0] p2_smul_37277_comb;
  wire [46:0] p2_smul_37280_comb;
  wire [46:0] p2_smul_37283_comb;
  wire [46:0] p2_smul_37286_comb;
  wire [31:0] p2_add_37471_comb;
  wire [31:0] p2_add_37472_comb;
  wire [31:0] p2_add_37473_comb;
  wire [31:0] p2_add_37474_comb;
  wire [31:0] p2_add_37475_comb;
  wire [31:0] p2_add_37476_comb;
  wire [31:0] p2_add_37477_comb;
  wire [31:0] p2_add_37478_comb;
  wire [31:0] p2_add_37479_comb;
  wire [31:0] p2_add_37480_comb;
  wire [31:0] p2_add_37481_comb;
  wire [31:0] p2_add_37482_comb;
  wire [31:0] p2_add_37483_comb;
  wire [31:0] p2_add_37484_comb;
  wire [31:0] p2_add_37485_comb;
  wire [31:0] p2_add_37486_comb;
  wire [15:0] p2_add_37535_comb;
  wire [15:0] p2_add_37536_comb;
  wire [15:0] p2_add_37537_comb;
  wire [15:0] p2_add_37538_comb;
  wire [15:0] p2_add_37539_comb;
  wire [15:0] p2_add_37540_comb;
  wire [15:0] p2_add_37541_comb;
  wire [15:0] p2_add_37542_comb;
  wire [15:0] p2_add_37543_comb;
  wire [15:0] p2_add_37544_comb;
  wire [15:0] p2_add_37545_comb;
  wire [15:0] p2_add_37546_comb;
  wire [15:0] p2_add_37547_comb;
  wire [15:0] p2_add_37548_comb;
  wire [15:0] p2_add_37549_comb;
  wire [15:0] p2_add_37550_comb;
  wire [15:0] p2_smul_37159_comb;
  wire [15:0] p2_sub_37160_comb;
  wire [15:0] p2_smul_37164_comb;
  wire [15:0] p2_sub_37165_comb;
  wire [15:0] p2_smul_37169_comb;
  wire [15:0] p2_sub_37170_comb;
  wire [15:0] p2_smul_37174_comb;
  wire [15:0] p2_sub_37175_comb;
  wire [15:0] p2_smul_37179_comb;
  wire [15:0] p2_sub_37180_comb;
  wire [15:0] p2_smul_37184_comb;
  wire [15:0] p2_sub_37185_comb;
  wire [15:0] p2_smul_37189_comb;
  wire [15:0] p2_sub_37190_comb;
  wire [15:0] p2_smul_37194_comb;
  wire [15:0] p2_sub_37195_comb;
  wire [15:0] p2_smul_37199_comb;
  wire [15:0] p2_sub_37200_comb;
  wire [15:0] p2_smul_37204_comb;
  wire [15:0] p2_sub_37205_comb;
  wire [15:0] p2_smul_37209_comb;
  wire [15:0] p2_sub_37210_comb;
  wire [15:0] p2_smul_37214_comb;
  wire [15:0] p2_sub_37215_comb;
  wire [15:0] p2_smul_37219_comb;
  wire [15:0] p2_sub_37220_comb;
  wire [15:0] p2_smul_37224_comb;
  wire [15:0] p2_sub_37225_comb;
  wire [15:0] p2_smul_37229_comb;
  wire [15:0] p2_sub_37230_comb;
  wire [15:0] p2_smul_37234_comb;
  wire [15:0] p2_sub_37235_comb;
  wire [15:0] p2_sub_37239_comb;
  wire [15:0] p2_sub_37242_comb;
  wire [15:0] p2_sub_37245_comb;
  wire [15:0] p2_sub_37248_comb;
  wire [15:0] p2_sub_37251_comb;
  wire [15:0] p2_sub_37254_comb;
  wire [15:0] p2_sub_37257_comb;
  wire [15:0] p2_sub_37260_comb;
  wire [15:0] p2_bit_slice_37263_comb;
  wire [15:0] p2_bit_slice_37266_comb;
  wire [15:0] p2_bit_slice_37269_comb;
  wire [15:0] p2_bit_slice_37272_comb;
  wire [15:0] p2_bit_slice_37275_comb;
  wire [15:0] p2_bit_slice_37278_comb;
  wire [15:0] p2_bit_slice_37281_comb;
  wire [15:0] p2_bit_slice_37284_comb;
  wire [15:0] p2_bit_slice_37287_comb;
  wire [15:0] p2_bit_slice_37289_comb;
  wire [15:0] p2_bit_slice_37291_comb;
  wire [15:0] p2_bit_slice_37293_comb;
  wire [15:0] p2_bit_slice_37295_comb;
  wire [15:0] p2_bit_slice_37297_comb;
  wire [15:0] p2_bit_slice_37299_comb;
  wire [15:0] p2_bit_slice_37301_comb;
  wire [15:0] p2_sub_37303_comb;
  wire [13:0] p2_bit_slice_37305_comb;
  wire [15:0] p2_sub_37306_comb;
  wire [13:0] p2_bit_slice_37308_comb;
  wire [15:0] p2_sub_37309_comb;
  wire [13:0] p2_bit_slice_37311_comb;
  wire [15:0] p2_sub_37312_comb;
  wire [13:0] p2_bit_slice_37314_comb;
  wire [15:0] p2_sub_37315_comb;
  wire [13:0] p2_bit_slice_37317_comb;
  wire [15:0] p2_sub_37318_comb;
  wire [13:0] p2_bit_slice_37320_comb;
  wire [15:0] p2_sub_37321_comb;
  wire [13:0] p2_bit_slice_37323_comb;
  wire [15:0] p2_sub_37324_comb;
  wire [13:0] p2_bit_slice_37326_comb;
  wire [15:0] p2_sub_37327_comb;
  wire [15:0] p2_sub_37329_comb;
  wire [15:0] p2_sub_37331_comb;
  wire [15:0] p2_sub_37333_comb;
  wire [15:0] p2_sub_37335_comb;
  wire [15:0] p2_sub_37337_comb;
  wire [15:0] p2_sub_37339_comb;
  wire [15:0] p2_sub_37341_comb;
  wire [15:0] p2_sub_37343_comb;
  wire [15:0] p2_sub_37344_comb;
  wire [15:0] p2_sub_37345_comb;
  wire [15:0] p2_sub_37346_comb;
  wire [15:0] p2_sub_37347_comb;
  wire [15:0] p2_sub_37348_comb;
  wire [15:0] p2_sub_37349_comb;
  wire [15:0] p2_sub_37350_comb;
  wire [15:0] p2_sub_37351_comb;
  wire [15:0] p2_sub_37352_comb;
  wire [15:0] p2_sub_37353_comb;
  wire [15:0] p2_sub_37354_comb;
  wire [15:0] p2_sub_37355_comb;
  wire [15:0] p2_sub_37356_comb;
  wire [15:0] p2_sub_37357_comb;
  wire [15:0] p2_sub_37358_comb;
  wire [15:0] p2_sub_37375_comb;
  wire [15:0] p2_sub_37376_comb;
  wire [15:0] p2_sub_37377_comb;
  wire [15:0] p2_sub_37378_comb;
  wire [15:0] p2_sub_37379_comb;
  wire [15:0] p2_sub_37380_comb;
  wire [15:0] p2_sub_37381_comb;
  wire [15:0] p2_sub_37382_comb;
  wire [15:0] p2_sub_37383_comb;
  wire [15:0] p2_sub_37384_comb;
  wire [15:0] p2_sub_37385_comb;
  wire [15:0] p2_sub_37386_comb;
  wire [15:0] p2_sub_37387_comb;
  wire [15:0] p2_sub_37388_comb;
  wire [15:0] p2_sub_37389_comb;
  wire [15:0] p2_sub_37390_comb;
  wire [15:0] p2_sub_37439_comb;
  wire [15:0] p2_sub_37441_comb;
  wire [15:0] p2_sub_37443_comb;
  wire [15:0] p2_sub_37445_comb;
  wire [15:0] p2_sub_37447_comb;
  wire [15:0] p2_sub_37449_comb;
  wire [15:0] p2_sub_37451_comb;
  wire [15:0] p2_sub_37453_comb;
  wire [15:0] p2_sub_37455_comb;
  wire [15:0] p2_sub_37457_comb;
  wire [15:0] p2_sub_37459_comb;
  wire [15:0] p2_sub_37461_comb;
  wire [15:0] p2_sub_37463_comb;
  wire [15:0] p2_sub_37465_comb;
  wire [15:0] p2_sub_37467_comb;
  wire [15:0] p2_sub_37469_comb;
  wire [15:0] p2_bit_slice_37487_comb;
  wire [15:0] p2_bit_slice_37488_comb;
  wire [15:0] p2_bit_slice_37489_comb;
  wire [15:0] p2_bit_slice_37490_comb;
  wire [15:0] p2_bit_slice_37491_comb;
  wire [15:0] p2_bit_slice_37492_comb;
  wire [15:0] p2_bit_slice_37493_comb;
  wire [15:0] p2_bit_slice_37494_comb;
  wire [15:0] p2_bit_slice_37495_comb;
  wire [15:0] p2_bit_slice_37496_comb;
  wire [15:0] p2_bit_slice_37497_comb;
  wire [15:0] p2_bit_slice_37498_comb;
  wire [15:0] p2_bit_slice_37499_comb;
  wire [15:0] p2_bit_slice_37500_comb;
  wire [15:0] p2_bit_slice_37501_comb;
  wire [15:0] p2_bit_slice_37502_comb;
  wire [15:0] p2_sub_37519_comb;
  wire [15:0] p2_sub_37520_comb;
  wire [15:0] p2_sub_37521_comb;
  wire [15:0] p2_sub_37522_comb;
  wire [15:0] p2_sub_37523_comb;
  wire [15:0] p2_sub_37524_comb;
  wire [15:0] p2_sub_37525_comb;
  wire [15:0] p2_sub_37526_comb;
  wire [15:0] p2_sub_37527_comb;
  wire [15:0] p2_sub_37528_comb;
  wire [15:0] p2_sub_37529_comb;
  wire [15:0] p2_sub_37530_comb;
  wire [15:0] p2_sub_37531_comb;
  wire [15:0] p2_sub_37532_comb;
  wire [15:0] p2_sub_37533_comb;
  wire [15:0] p2_sub_37534_comb;
  wire [15:0] p2_add_37551_comb;
  wire [15:0] p2_add_37552_comb;
  wire [15:0] p2_add_37553_comb;
  wire [15:0] p2_add_37554_comb;
  wire [15:0] p2_add_37555_comb;
  wire [15:0] p2_add_37556_comb;
  wire [15:0] p2_add_37557_comb;
  wire [15:0] p2_add_37558_comb;
  wire [15:0] p2_add_37559_comb;
  wire [15:0] p2_add_37560_comb;
  wire [15:0] p2_add_37561_comb;
  wire [15:0] p2_add_37562_comb;
  wire [15:0] p2_add_37563_comb;
  wire [15:0] p2_add_37564_comb;
  wire [15:0] p2_add_37565_comb;
  wire [15:0] p2_add_37566_comb;
  wire [15:0] p2_add_37567_comb;
  wire [15:0] p2_add_37568_comb;
  wire [15:0] p2_add_37569_comb;
  wire [15:0] p2_add_37570_comb;
  wire [15:0] p2_add_37571_comb;
  wire [15:0] p2_add_37572_comb;
  wire [15:0] p2_add_37573_comb;
  wire [15:0] p2_add_37574_comb;
  assign p2_sign_ext_36615_comb = {{16{p1_neg_36551[15]}}, p1_neg_36551};
  assign p2_sign_ext_36616_comb = {{16{p1_neg_36552[15]}}, p1_neg_36552};
  assign p2_sign_ext_36617_comb = {{16{p1_neg_36553[15]}}, p1_neg_36553};
  assign p2_sign_ext_36618_comb = {{16{p1_neg_36554[15]}}, p1_neg_36554};
  assign p2_sign_ext_36619_comb = {{16{p1_neg_36555[15]}}, p1_neg_36555};
  assign p2_sign_ext_36620_comb = {{16{p1_neg_36556[15]}}, p1_neg_36556};
  assign p2_sign_ext_36621_comb = {{16{p1_neg_36557[15]}}, p1_neg_36557};
  assign p2_sign_ext_36622_comb = {{16{p1_neg_36558[15]}}, p1_neg_36558};
  assign p2_add_36687_comb = p1_sign_ext_36559 + {31'h0000_0000, p1_sign_ext_36559[31]};
  assign p2_smul_33601_NarrowedMult__comb = smul47b_16b_x_31b(p1_neg_36543, 31'h2aaa_aaab);
  assign p2_add_36692_comb = p1_sign_ext_36560 + {31'h0000_0000, p1_sign_ext_36560[31]};
  assign p2_smul_33603_NarrowedMult__comb = smul47b_16b_x_31b(p1_neg_36544, 31'h2aaa_aaab);
  assign p2_add_36697_comb = p1_sign_ext_36561 + {31'h0000_0000, p1_sign_ext_36561[31]};
  assign p2_smul_33605_NarrowedMult__comb = smul47b_16b_x_31b(p1_neg_36545, 31'h2aaa_aaab);
  assign p2_add_36702_comb = p1_sign_ext_36562 + {31'h0000_0000, p1_sign_ext_36562[31]};
  assign p2_smul_33607_NarrowedMult__comb = smul47b_16b_x_31b(p1_neg_36546, 31'h2aaa_aaab);
  assign p2_add_36707_comb = p1_sign_ext_36563 + {31'h0000_0000, p1_sign_ext_36563[31]};
  assign p2_smul_33609_NarrowedMult__comb = smul47b_16b_x_31b(p1_neg_36547, 31'h2aaa_aaab);
  assign p2_add_36712_comb = p1_sign_ext_36564 + {31'h0000_0000, p1_sign_ext_36564[31]};
  assign p2_smul_33611_NarrowedMult__comb = smul47b_16b_x_31b(p1_neg_36548, 31'h2aaa_aaab);
  assign p2_add_36717_comb = p1_sign_ext_36565 + {31'h0000_0000, p1_sign_ext_36565[31]};
  assign p2_smul_33613_NarrowedMult__comb = smul47b_16b_x_31b(p1_neg_36549, 31'h2aaa_aaab);
  assign p2_add_36722_comb = p1_sign_ext_36566 + {31'h0000_0000, p1_sign_ext_36566[31]};
  assign p2_smul_33615_NarrowedMult__comb = smul47b_16b_x_31b(p1_neg_36550, 31'h2aaa_aaab);
  assign p2_add_36727_comb = p2_sign_ext_36615_comb + {31'h0000_0000, p2_sign_ext_36615_comb[31]};
  assign p2_smul_33617_NarrowedMult__comb = smul47b_16b_x_31b(p1_neg_36551, 31'h2aaa_aaab);
  assign p2_add_36732_comb = p2_sign_ext_36616_comb + {31'h0000_0000, p2_sign_ext_36616_comb[31]};
  assign p2_smul_33619_NarrowedMult__comb = smul47b_16b_x_31b(p1_neg_36552, 31'h2aaa_aaab);
  assign p2_add_36737_comb = p2_sign_ext_36617_comb + {31'h0000_0000, p2_sign_ext_36617_comb[31]};
  assign p2_smul_33621_NarrowedMult__comb = smul47b_16b_x_31b(p1_neg_36553, 31'h2aaa_aaab);
  assign p2_add_36742_comb = p2_sign_ext_36618_comb + {31'h0000_0000, p2_sign_ext_36618_comb[31]};
  assign p2_smul_33623_NarrowedMult__comb = smul47b_16b_x_31b(p1_neg_36554, 31'h2aaa_aaab);
  assign p2_add_36747_comb = p2_sign_ext_36619_comb + {31'h0000_0000, p2_sign_ext_36619_comb[31]};
  assign p2_smul_33625_NarrowedMult__comb = smul47b_16b_x_31b(p1_neg_36555, 31'h2aaa_aaab);
  assign p2_add_36752_comb = p2_sign_ext_36620_comb + {31'h0000_0000, p2_sign_ext_36620_comb[31]};
  assign p2_smul_33627_NarrowedMult__comb = smul47b_16b_x_31b(p1_neg_36556, 31'h2aaa_aaab);
  assign p2_add_36757_comb = p2_sign_ext_36621_comb + {31'h0000_0000, p2_sign_ext_36621_comb[31]};
  assign p2_smul_33629_NarrowedMult__comb = smul47b_16b_x_31b(p1_neg_36557, 31'h2aaa_aaab);
  assign p2_add_36762_comb = p2_sign_ext_36622_comb + {31'h0000_0000, p2_sign_ext_36622_comb[31]};
  assign p2_smul_33631_NarrowedMult__comb = smul47b_16b_x_31b(p1_neg_36558, 31'h2aaa_aaab);
  assign p2_sign_ext_36769_comb = {16{p1_sign_ext_36559[31]}};
  assign p2_smul_36771_comb = smul48b_16b_x_32b(p1_neg_36543, 32'h6666_6667);
  assign p2_sign_ext_36774_comb = {16{p1_sign_ext_36560[31]}};
  assign p2_smul_36776_comb = smul48b_16b_x_32b(p1_neg_36544, 32'h6666_6667);
  assign p2_sign_ext_36779_comb = {16{p1_sign_ext_36561[31]}};
  assign p2_smul_36781_comb = smul48b_16b_x_32b(p1_neg_36545, 32'h6666_6667);
  assign p2_sign_ext_36784_comb = {16{p1_sign_ext_36562[31]}};
  assign p2_smul_36786_comb = smul48b_16b_x_32b(p1_neg_36546, 32'h6666_6667);
  assign p2_sign_ext_36789_comb = {16{p1_sign_ext_36563[31]}};
  assign p2_smul_36791_comb = smul48b_16b_x_32b(p1_neg_36547, 32'h6666_6667);
  assign p2_sign_ext_36794_comb = {16{p1_sign_ext_36564[31]}};
  assign p2_smul_36796_comb = smul48b_16b_x_32b(p1_neg_36548, 32'h6666_6667);
  assign p2_sign_ext_36799_comb = {16{p1_sign_ext_36565[31]}};
  assign p2_smul_36801_comb = smul48b_16b_x_32b(p1_neg_36549, 32'h6666_6667);
  assign p2_sign_ext_36804_comb = {16{p1_sign_ext_36566[31]}};
  assign p2_smul_36806_comb = smul48b_16b_x_32b(p1_neg_36550, 32'h6666_6667);
  assign p2_sign_ext_36809_comb = {16{p2_sign_ext_36615_comb[31]}};
  assign p2_smul_36811_comb = smul48b_16b_x_32b(p1_neg_36551, 32'h6666_6667);
  assign p2_sign_ext_36814_comb = {16{p2_sign_ext_36616_comb[31]}};
  assign p2_smul_36816_comb = smul48b_16b_x_32b(p1_neg_36552, 32'h6666_6667);
  assign p2_sign_ext_36819_comb = {16{p2_sign_ext_36617_comb[31]}};
  assign p2_smul_36821_comb = smul48b_16b_x_32b(p1_neg_36553, 32'h6666_6667);
  assign p2_sign_ext_36824_comb = {16{p2_sign_ext_36618_comb[31]}};
  assign p2_smul_36826_comb = smul48b_16b_x_32b(p1_neg_36554, 32'h6666_6667);
  assign p2_sign_ext_36829_comb = {16{p2_sign_ext_36619_comb[31]}};
  assign p2_smul_36831_comb = smul48b_16b_x_32b(p1_neg_36555, 32'h6666_6667);
  assign p2_sign_ext_36834_comb = {16{p2_sign_ext_36620_comb[31]}};
  assign p2_smul_36836_comb = smul48b_16b_x_32b(p1_neg_36556, 32'h6666_6667);
  assign p2_sign_ext_36839_comb = {16{p2_sign_ext_36621_comb[31]}};
  assign p2_smul_36841_comb = smul48b_16b_x_32b(p1_neg_36557, 32'h6666_6667);
  assign p2_sign_ext_36844_comb = {16{p2_sign_ext_36622_comb[31]}};
  assign p2_smul_36846_comb = smul48b_16b_x_32b(p1_neg_36558, 32'h6666_6667);
  assign p2_smul_36847_comb = smul16b_16b_x_16b(p1_neg_36543, p2_add_36687_comb[16:1]);
  assign p2_sub_36848_comb = p2_smul_33601_NarrowedMult__comb[46:31] - p2_sign_ext_36769_comb;
  assign p2_add_36849_comb = p1_sign_ext_36559 + {30'h0000_0000, {2{p1_sign_ext_36559[31]}}};
  assign p2_sign_ext_36850_comb = {{16{p2_smul_36771_comb[47]}}, p2_smul_36771_comb};
  assign p2_smul_36852_comb = smul16b_16b_x_16b(p1_neg_36544, p2_add_36692_comb[16:1]);
  assign p2_sub_36853_comb = p2_smul_33603_NarrowedMult__comb[46:31] - p2_sign_ext_36774_comb;
  assign p2_add_36854_comb = p1_sign_ext_36560 + {30'h0000_0000, {2{p1_sign_ext_36560[31]}}};
  assign p2_sign_ext_36855_comb = {{16{p2_smul_36776_comb[47]}}, p2_smul_36776_comb};
  assign p2_smul_36857_comb = smul16b_16b_x_16b(p1_neg_36545, p2_add_36697_comb[16:1]);
  assign p2_sub_36858_comb = p2_smul_33605_NarrowedMult__comb[46:31] - p2_sign_ext_36779_comb;
  assign p2_add_36859_comb = p1_sign_ext_36561 + {30'h0000_0000, {2{p1_sign_ext_36561[31]}}};
  assign p2_sign_ext_36860_comb = {{16{p2_smul_36781_comb[47]}}, p2_smul_36781_comb};
  assign p2_smul_36862_comb = smul16b_16b_x_16b(p1_neg_36546, p2_add_36702_comb[16:1]);
  assign p2_sub_36863_comb = p2_smul_33607_NarrowedMult__comb[46:31] - p2_sign_ext_36784_comb;
  assign p2_add_36864_comb = p1_sign_ext_36562 + {30'h0000_0000, {2{p1_sign_ext_36562[31]}}};
  assign p2_sign_ext_36865_comb = {{16{p2_smul_36786_comb[47]}}, p2_smul_36786_comb};
  assign p2_smul_36867_comb = smul16b_16b_x_16b(p1_neg_36547, p2_add_36707_comb[16:1]);
  assign p2_sub_36868_comb = p2_smul_33609_NarrowedMult__comb[46:31] - p2_sign_ext_36789_comb;
  assign p2_add_36869_comb = p1_sign_ext_36563 + {30'h0000_0000, {2{p1_sign_ext_36563[31]}}};
  assign p2_sign_ext_36870_comb = {{16{p2_smul_36791_comb[47]}}, p2_smul_36791_comb};
  assign p2_smul_36872_comb = smul16b_16b_x_16b(p1_neg_36548, p2_add_36712_comb[16:1]);
  assign p2_sub_36873_comb = p2_smul_33611_NarrowedMult__comb[46:31] - p2_sign_ext_36794_comb;
  assign p2_add_36874_comb = p1_sign_ext_36564 + {30'h0000_0000, {2{p1_sign_ext_36564[31]}}};
  assign p2_sign_ext_36875_comb = {{16{p2_smul_36796_comb[47]}}, p2_smul_36796_comb};
  assign p2_smul_36877_comb = smul16b_16b_x_16b(p1_neg_36549, p2_add_36717_comb[16:1]);
  assign p2_sub_36878_comb = p2_smul_33613_NarrowedMult__comb[46:31] - p2_sign_ext_36799_comb;
  assign p2_add_36879_comb = p1_sign_ext_36565 + {30'h0000_0000, {2{p1_sign_ext_36565[31]}}};
  assign p2_sign_ext_36880_comb = {{16{p2_smul_36801_comb[47]}}, p2_smul_36801_comb};
  assign p2_smul_36882_comb = smul16b_16b_x_16b(p1_neg_36550, p2_add_36722_comb[16:1]);
  assign p2_sub_36883_comb = p2_smul_33615_NarrowedMult__comb[46:31] - p2_sign_ext_36804_comb;
  assign p2_add_36884_comb = p1_sign_ext_36566 + {30'h0000_0000, {2{p1_sign_ext_36566[31]}}};
  assign p2_sign_ext_36885_comb = {{16{p2_smul_36806_comb[47]}}, p2_smul_36806_comb};
  assign p2_smul_36887_comb = smul16b_16b_x_16b(p1_neg_36551, p2_add_36727_comb[16:1]);
  assign p2_sub_36888_comb = p2_smul_33617_NarrowedMult__comb[46:31] - p2_sign_ext_36809_comb;
  assign p2_add_36889_comb = p2_sign_ext_36615_comb + {30'h0000_0000, {2{p2_sign_ext_36615_comb[31]}}};
  assign p2_sign_ext_36890_comb = {{16{p2_smul_36811_comb[47]}}, p2_smul_36811_comb};
  assign p2_smul_36892_comb = smul16b_16b_x_16b(p1_neg_36552, p2_add_36732_comb[16:1]);
  assign p2_sub_36893_comb = p2_smul_33619_NarrowedMult__comb[46:31] - p2_sign_ext_36814_comb;
  assign p2_add_36894_comb = p2_sign_ext_36616_comb + {30'h0000_0000, {2{p2_sign_ext_36616_comb[31]}}};
  assign p2_sign_ext_36895_comb = {{16{p2_smul_36816_comb[47]}}, p2_smul_36816_comb};
  assign p2_smul_36897_comb = smul16b_16b_x_16b(p1_neg_36553, p2_add_36737_comb[16:1]);
  assign p2_sub_36898_comb = p2_smul_33621_NarrowedMult__comb[46:31] - p2_sign_ext_36819_comb;
  assign p2_add_36899_comb = p2_sign_ext_36617_comb + {30'h0000_0000, {2{p2_sign_ext_36617_comb[31]}}};
  assign p2_sign_ext_36900_comb = {{16{p2_smul_36821_comb[47]}}, p2_smul_36821_comb};
  assign p2_smul_36902_comb = smul16b_16b_x_16b(p1_neg_36554, p2_add_36742_comb[16:1]);
  assign p2_sub_36903_comb = p2_smul_33623_NarrowedMult__comb[46:31] - p2_sign_ext_36824_comb;
  assign p2_add_36904_comb = p2_sign_ext_36618_comb + {30'h0000_0000, {2{p2_sign_ext_36618_comb[31]}}};
  assign p2_sign_ext_36905_comb = {{16{p2_smul_36826_comb[47]}}, p2_smul_36826_comb};
  assign p2_smul_36907_comb = smul16b_16b_x_16b(p1_neg_36555, p2_add_36747_comb[16:1]);
  assign p2_sub_36908_comb = p2_smul_33625_NarrowedMult__comb[46:31] - p2_sign_ext_36829_comb;
  assign p2_add_36909_comb = p2_sign_ext_36619_comb + {30'h0000_0000, {2{p2_sign_ext_36619_comb[31]}}};
  assign p2_sign_ext_36910_comb = {{16{p2_smul_36831_comb[47]}}, p2_smul_36831_comb};
  assign p2_smul_36912_comb = smul16b_16b_x_16b(p1_neg_36556, p2_add_36752_comb[16:1]);
  assign p2_sub_36913_comb = p2_smul_33627_NarrowedMult__comb[46:31] - p2_sign_ext_36834_comb;
  assign p2_add_36914_comb = p2_sign_ext_36620_comb + {30'h0000_0000, {2{p2_sign_ext_36620_comb[31]}}};
  assign p2_sign_ext_36915_comb = {{16{p2_smul_36836_comb[47]}}, p2_smul_36836_comb};
  assign p2_smul_36917_comb = smul16b_16b_x_16b(p1_neg_36557, p2_add_36757_comb[16:1]);
  assign p2_sub_36918_comb = p2_smul_33629_NarrowedMult__comb[46:31] - p2_sign_ext_36839_comb;
  assign p2_add_36919_comb = p2_sign_ext_36621_comb + {30'h0000_0000, {2{p2_sign_ext_36621_comb[31]}}};
  assign p2_sign_ext_36920_comb = {{16{p2_smul_36841_comb[47]}}, p2_smul_36841_comb};
  assign p2_smul_36922_comb = smul16b_16b_x_16b(p1_neg_36558, p2_add_36762_comb[16:1]);
  assign p2_sub_36923_comb = p2_smul_33631_NarrowedMult__comb[46:31] - p2_sign_ext_36844_comb;
  assign p2_add_36924_comb = p2_sign_ext_36622_comb + {30'h0000_0000, {2{p2_sign_ext_36622_comb[31]}}};
  assign p2_sign_ext_36925_comb = {{16{p2_smul_36846_comb[47]}}, p2_smul_36846_comb};
  assign p2_smul_36927_comb = smul16b_16b_x_16b(p2_smul_36847_comb, p2_sub_36848_comb);
  assign p2_sign_ext_36930_comb = {{16{p2_smul_33601_NarrowedMult__comb[46]}}, p2_smul_33601_NarrowedMult__comb};
  assign p2_smul_36931_comb = smul49b_16b_x_33b(p1_neg_36543, 33'h0_9249_2493);
  assign p2_smul_36932_comb = smul16b_16b_x_16b(p2_smul_36852_comb, p2_sub_36853_comb);
  assign p2_sign_ext_36935_comb = {{16{p2_smul_33603_NarrowedMult__comb[46]}}, p2_smul_33603_NarrowedMult__comb};
  assign p2_smul_36936_comb = smul49b_16b_x_33b(p1_neg_36544, 33'h0_9249_2493);
  assign p2_smul_36937_comb = smul16b_16b_x_16b(p2_smul_36857_comb, p2_sub_36858_comb);
  assign p2_sign_ext_36940_comb = {{16{p2_smul_33605_NarrowedMult__comb[46]}}, p2_smul_33605_NarrowedMult__comb};
  assign p2_smul_36941_comb = smul49b_16b_x_33b(p1_neg_36545, 33'h0_9249_2493);
  assign p2_smul_36942_comb = smul16b_16b_x_16b(p2_smul_36862_comb, p2_sub_36863_comb);
  assign p2_sign_ext_36945_comb = {{16{p2_smul_33607_NarrowedMult__comb[46]}}, p2_smul_33607_NarrowedMult__comb};
  assign p2_smul_36946_comb = smul49b_16b_x_33b(p1_neg_36546, 33'h0_9249_2493);
  assign p2_smul_36947_comb = smul16b_16b_x_16b(p2_smul_36867_comb, p2_sub_36868_comb);
  assign p2_sign_ext_36950_comb = {{16{p2_smul_33609_NarrowedMult__comb[46]}}, p2_smul_33609_NarrowedMult__comb};
  assign p2_smul_36951_comb = smul49b_16b_x_33b(p1_neg_36547, 33'h0_9249_2493);
  assign p2_smul_36952_comb = smul16b_16b_x_16b(p2_smul_36872_comb, p2_sub_36873_comb);
  assign p2_sign_ext_36955_comb = {{16{p2_smul_33611_NarrowedMult__comb[46]}}, p2_smul_33611_NarrowedMult__comb};
  assign p2_smul_36956_comb = smul49b_16b_x_33b(p1_neg_36548, 33'h0_9249_2493);
  assign p2_smul_36957_comb = smul16b_16b_x_16b(p2_smul_36877_comb, p2_sub_36878_comb);
  assign p2_sign_ext_36960_comb = {{16{p2_smul_33613_NarrowedMult__comb[46]}}, p2_smul_33613_NarrowedMult__comb};
  assign p2_smul_36961_comb = smul49b_16b_x_33b(p1_neg_36549, 33'h0_9249_2493);
  assign p2_smul_36962_comb = smul16b_16b_x_16b(p2_smul_36882_comb, p2_sub_36883_comb);
  assign p2_sign_ext_36965_comb = {{16{p2_smul_33615_NarrowedMult__comb[46]}}, p2_smul_33615_NarrowedMult__comb};
  assign p2_smul_36966_comb = smul49b_16b_x_33b(p1_neg_36550, 33'h0_9249_2493);
  assign p2_smul_36971_comb = smul49b_16b_x_33b(p1_neg_36551, 33'h0_9249_2493);
  assign p2_smul_36976_comb = smul49b_16b_x_33b(p1_neg_36552, 33'h0_9249_2493);
  assign p2_smul_36981_comb = smul49b_16b_x_33b(p1_neg_36553, 33'h0_9249_2493);
  assign p2_smul_36986_comb = smul49b_16b_x_33b(p1_neg_36554, 33'h0_9249_2493);
  assign p2_smul_36991_comb = smul49b_16b_x_33b(p1_neg_36555, 33'h0_9249_2493);
  assign p2_smul_36996_comb = smul49b_16b_x_33b(p1_neg_36556, 33'h0_9249_2493);
  assign p2_smul_37001_comb = smul49b_16b_x_33b(p1_neg_36557, 33'h0_9249_2493);
  assign p2_smul_37006_comb = smul49b_16b_x_33b(p1_neg_36558, 33'h0_9249_2493);
  assign p2_smul_37123_comb = smul47b_16b_x_31b(p1_neg_36543, 31'h38e3_8e39);
  assign p2_smul_37128_comb = smul47b_16b_x_31b(p1_neg_36544, 31'h38e3_8e39);
  assign p2_smul_37133_comb = smul47b_16b_x_31b(p1_neg_36545, 31'h38e3_8e39);
  assign p2_smul_37138_comb = smul47b_16b_x_31b(p1_neg_36546, 31'h38e3_8e39);
  assign p2_smul_37143_comb = smul47b_16b_x_31b(p1_neg_36547, 31'h38e3_8e39);
  assign p2_smul_37148_comb = smul47b_16b_x_31b(p1_neg_36548, 31'h38e3_8e39);
  assign p2_smul_37153_comb = smul47b_16b_x_31b(p1_neg_36549, 31'h38e3_8e39);
  assign p2_smul_37158_comb = smul47b_16b_x_31b(p1_neg_36550, 31'h38e3_8e39);
  assign p2_smul_37163_comb = smul47b_16b_x_31b(p1_neg_36551, 31'h38e3_8e39);
  assign p2_smul_37168_comb = smul47b_16b_x_31b(p1_neg_36552, 31'h38e3_8e39);
  assign p2_smul_37173_comb = smul47b_16b_x_31b(p1_neg_36553, 31'h38e3_8e39);
  assign p2_smul_37178_comb = smul47b_16b_x_31b(p1_neg_36554, 31'h38e3_8e39);
  assign p2_smul_37183_comb = smul47b_16b_x_31b(p1_neg_36555, 31'h38e3_8e39);
  assign p2_smul_37188_comb = smul47b_16b_x_31b(p1_neg_36556, 31'h38e3_8e39);
  assign p2_smul_37193_comb = smul47b_16b_x_31b(p1_neg_36557, 31'h38e3_8e39);
  assign p2_smul_37198_comb = smul47b_16b_x_31b(p1_neg_36558, 31'h38e3_8e39);
  assign p2_smul_36967_comb = smul16b_16b_x_16b(p2_smul_36887_comb, p2_sub_36888_comb);
  assign p2_sign_ext_36970_comb = {{16{p2_smul_33617_NarrowedMult__comb[46]}}, p2_smul_33617_NarrowedMult__comb};
  assign p2_smul_36972_comb = smul16b_16b_x_16b(p2_smul_36892_comb, p2_sub_36893_comb);
  assign p2_sign_ext_36975_comb = {{16{p2_smul_33619_NarrowedMult__comb[46]}}, p2_smul_33619_NarrowedMult__comb};
  assign p2_smul_36977_comb = smul16b_16b_x_16b(p2_smul_36897_comb, p2_sub_36898_comb);
  assign p2_sign_ext_36980_comb = {{16{p2_smul_33621_NarrowedMult__comb[46]}}, p2_smul_33621_NarrowedMult__comb};
  assign p2_smul_36982_comb = smul16b_16b_x_16b(p2_smul_36902_comb, p2_sub_36903_comb);
  assign p2_sign_ext_36985_comb = {{16{p2_smul_33623_NarrowedMult__comb[46]}}, p2_smul_33623_NarrowedMult__comb};
  assign p2_smul_36987_comb = smul16b_16b_x_16b(p2_smul_36907_comb, p2_sub_36908_comb);
  assign p2_sign_ext_36990_comb = {{16{p2_smul_33625_NarrowedMult__comb[46]}}, p2_smul_33625_NarrowedMult__comb};
  assign p2_smul_36992_comb = smul16b_16b_x_16b(p2_smul_36912_comb, p2_sub_36913_comb);
  assign p2_sign_ext_36995_comb = {{16{p2_smul_33627_NarrowedMult__comb[46]}}, p2_smul_33627_NarrowedMult__comb};
  assign p2_smul_36997_comb = smul16b_16b_x_16b(p2_smul_36917_comb, p2_sub_36918_comb);
  assign p2_sign_ext_37000_comb = {{16{p2_smul_33629_NarrowedMult__comb[46]}}, p2_smul_33629_NarrowedMult__comb};
  assign p2_smul_37002_comb = smul16b_16b_x_16b(p2_smul_36922_comb, p2_sub_36923_comb);
  assign p2_sign_ext_37005_comb = {{16{p2_smul_33631_NarrowedMult__comb[46]}}, p2_smul_33631_NarrowedMult__comb};
  assign p2_smul_37007_comb = smul16b_16b_x_16b(p2_smul_36927_comb, p2_add_36849_comb[17:2]);
  assign p2_sub_37008_comb = p2_sign_ext_36850_comb[48:33] - p2_sign_ext_36769_comb;
  assign p2_sign_ext_37010_comb = {{16{p2_smul_36931_comb[48]}}, p2_smul_36931_comb};
  assign p2_smul_37014_comb = smul16b_16b_x_16b(p2_smul_36932_comb, p2_add_36854_comb[17:2]);
  assign p2_sub_37015_comb = p2_sign_ext_36855_comb[48:33] - p2_sign_ext_36774_comb;
  assign p2_sign_ext_37017_comb = {{16{p2_smul_36936_comb[48]}}, p2_smul_36936_comb};
  assign p2_smul_37021_comb = smul16b_16b_x_16b(p2_smul_36937_comb, p2_add_36859_comb[17:2]);
  assign p2_sub_37022_comb = p2_sign_ext_36860_comb[48:33] - p2_sign_ext_36779_comb;
  assign p2_sign_ext_37024_comb = {{16{p2_smul_36941_comb[48]}}, p2_smul_36941_comb};
  assign p2_smul_37028_comb = smul16b_16b_x_16b(p2_smul_36942_comb, p2_add_36864_comb[17:2]);
  assign p2_sub_37029_comb = p2_sign_ext_36865_comb[48:33] - p2_sign_ext_36784_comb;
  assign p2_sign_ext_37031_comb = {{16{p2_smul_36946_comb[48]}}, p2_smul_36946_comb};
  assign p2_smul_37035_comb = smul16b_16b_x_16b(p2_smul_36947_comb, p2_add_36869_comb[17:2]);
  assign p2_sub_37036_comb = p2_sign_ext_36870_comb[48:33] - p2_sign_ext_36789_comb;
  assign p2_sign_ext_37038_comb = {{16{p2_smul_36951_comb[48]}}, p2_smul_36951_comb};
  assign p2_smul_37042_comb = smul16b_16b_x_16b(p2_smul_36952_comb, p2_add_36874_comb[17:2]);
  assign p2_sub_37043_comb = p2_sign_ext_36875_comb[48:33] - p2_sign_ext_36794_comb;
  assign p2_sign_ext_37045_comb = {{16{p2_smul_36956_comb[48]}}, p2_smul_36956_comb};
  assign p2_smul_37049_comb = smul16b_16b_x_16b(p2_smul_36957_comb, p2_add_36879_comb[17:2]);
  assign p2_sub_37050_comb = p2_sign_ext_36880_comb[48:33] - p2_sign_ext_36799_comb;
  assign p2_sign_ext_37052_comb = {{16{p2_smul_36961_comb[48]}}, p2_smul_36961_comb};
  assign p2_smul_37056_comb = smul16b_16b_x_16b(p2_smul_36962_comb, p2_add_36884_comb[17:2]);
  assign p2_sub_37057_comb = p2_sign_ext_36885_comb[48:33] - p2_sign_ext_36804_comb;
  assign p2_sign_ext_37059_comb = {{16{p2_smul_36966_comb[48]}}, p2_smul_36966_comb};
  assign p2_sign_ext_37066_comb = {{16{p2_smul_36971_comb[48]}}, p2_smul_36971_comb};
  assign p2_sign_ext_37073_comb = {{16{p2_smul_36976_comb[48]}}, p2_smul_36976_comb};
  assign p2_sign_ext_37080_comb = {{16{p2_smul_36981_comb[48]}}, p2_smul_36981_comb};
  assign p2_sign_ext_37087_comb = {{16{p2_smul_36986_comb[48]}}, p2_smul_36986_comb};
  assign p2_sign_ext_37094_comb = {{16{p2_smul_36991_comb[48]}}, p2_smul_36991_comb};
  assign p2_sign_ext_37101_comb = {{16{p2_smul_36996_comb[48]}}, p2_smul_36996_comb};
  assign p2_sign_ext_37108_comb = {{16{p2_smul_37001_comb[48]}}, p2_smul_37001_comb};
  assign p2_sign_ext_37115_comb = {{16{p2_smul_37006_comb[48]}}, p2_smul_37006_comb};
  assign p2_sign_ext_37202_comb = {{16{p2_smul_37123_comb[46]}}, p2_smul_37123_comb};
  assign p2_sign_ext_37207_comb = {{16{p2_smul_37128_comb[46]}}, p2_smul_37128_comb};
  assign p2_sign_ext_37212_comb = {{16{p2_smul_37133_comb[46]}}, p2_smul_37133_comb};
  assign p2_sign_ext_37217_comb = {{16{p2_smul_37138_comb[46]}}, p2_smul_37138_comb};
  assign p2_sign_ext_37222_comb = {{16{p2_smul_37143_comb[46]}}, p2_smul_37143_comb};
  assign p2_sign_ext_37227_comb = {{16{p2_smul_37148_comb[46]}}, p2_smul_37148_comb};
  assign p2_sign_ext_37232_comb = {{16{p2_smul_37153_comb[46]}}, p2_smul_37153_comb};
  assign p2_sign_ext_37237_comb = {{16{p2_smul_37158_comb[46]}}, p2_smul_37158_comb};
  assign p2_sign_ext_37241_comb = {{16{p2_smul_37163_comb[46]}}, p2_smul_37163_comb};
  assign p2_sign_ext_37244_comb = {{16{p2_smul_37168_comb[46]}}, p2_smul_37168_comb};
  assign p2_sign_ext_37247_comb = {{16{p2_smul_37173_comb[46]}}, p2_smul_37173_comb};
  assign p2_sign_ext_37250_comb = {{16{p2_smul_37178_comb[46]}}, p2_smul_37178_comb};
  assign p2_sign_ext_37253_comb = {{16{p2_smul_37183_comb[46]}}, p2_smul_37183_comb};
  assign p2_sign_ext_37256_comb = {{16{p2_smul_37188_comb[46]}}, p2_smul_37188_comb};
  assign p2_sign_ext_37259_comb = {{16{p2_smul_37193_comb[46]}}, p2_smul_37193_comb};
  assign p2_sign_ext_37262_comb = {{16{p2_smul_37198_comb[46]}}, p2_smul_37198_comb};
  assign p2_smul_37063_comb = smul16b_16b_x_16b(p2_smul_36967_comb, p2_add_36889_comb[17:2]);
  assign p2_sub_37064_comb = p2_sign_ext_36890_comb[48:33] - p2_sign_ext_36809_comb;
  assign p2_smul_37070_comb = smul16b_16b_x_16b(p2_smul_36972_comb, p2_add_36894_comb[17:2]);
  assign p2_sub_37071_comb = p2_sign_ext_36895_comb[48:33] - p2_sign_ext_36814_comb;
  assign p2_smul_37077_comb = smul16b_16b_x_16b(p2_smul_36977_comb, p2_add_36899_comb[17:2]);
  assign p2_sub_37078_comb = p2_sign_ext_36900_comb[48:33] - p2_sign_ext_36819_comb;
  assign p2_smul_37084_comb = smul16b_16b_x_16b(p2_smul_36982_comb, p2_add_36904_comb[17:2]);
  assign p2_sub_37085_comb = p2_sign_ext_36905_comb[48:33] - p2_sign_ext_36824_comb;
  assign p2_smul_37091_comb = smul16b_16b_x_16b(p2_smul_36987_comb, p2_add_36909_comb[17:2]);
  assign p2_sub_37092_comb = p2_sign_ext_36910_comb[48:33] - p2_sign_ext_36829_comb;
  assign p2_smul_37098_comb = smul16b_16b_x_16b(p2_smul_36992_comb, p2_add_36914_comb[17:2]);
  assign p2_sub_37099_comb = p2_sign_ext_36915_comb[48:33] - p2_sign_ext_36834_comb;
  assign p2_smul_37105_comb = smul16b_16b_x_16b(p2_smul_36997_comb, p2_add_36919_comb[17:2]);
  assign p2_sub_37106_comb = p2_sign_ext_36920_comb[48:33] - p2_sign_ext_36839_comb;
  assign p2_smul_37112_comb = smul16b_16b_x_16b(p2_smul_37002_comb, p2_add_36924_comb[17:2]);
  assign p2_sub_37113_comb = p2_sign_ext_36925_comb[48:33] - p2_sign_ext_36844_comb;
  assign p2_smul_37119_comb = smul16b_16b_x_16b(p2_smul_37007_comb, p2_sub_37008_comb);
  assign p2_sub_37120_comb = p2_sign_ext_36930_comb[47:32] - p2_sign_ext_36769_comb;
  assign p2_smul_37124_comb = smul16b_16b_x_16b(p2_smul_37014_comb, p2_sub_37015_comb);
  assign p2_sub_37125_comb = p2_sign_ext_36935_comb[47:32] - p2_sign_ext_36774_comb;
  assign p2_smul_37129_comb = smul16b_16b_x_16b(p2_smul_37021_comb, p2_sub_37022_comb);
  assign p2_sub_37130_comb = p2_sign_ext_36940_comb[47:32] - p2_sign_ext_36779_comb;
  assign p2_smul_37134_comb = smul16b_16b_x_16b(p2_smul_37028_comb, p2_sub_37029_comb);
  assign p2_sub_37135_comb = p2_sign_ext_36945_comb[47:32] - p2_sign_ext_36784_comb;
  assign p2_smul_37139_comb = smul16b_16b_x_16b(p2_smul_37035_comb, p2_sub_37036_comb);
  assign p2_sub_37140_comb = p2_sign_ext_36950_comb[47:32] - p2_sign_ext_36789_comb;
  assign p2_smul_37144_comb = smul16b_16b_x_16b(p2_smul_37042_comb, p2_sub_37043_comb);
  assign p2_sub_37145_comb = p2_sign_ext_36955_comb[47:32] - p2_sign_ext_36794_comb;
  assign p2_smul_37149_comb = smul16b_16b_x_16b(p2_smul_37049_comb, p2_sub_37050_comb);
  assign p2_sub_37150_comb = p2_sign_ext_36960_comb[47:32] - p2_sign_ext_36799_comb;
  assign p2_smul_37154_comb = smul16b_16b_x_16b(p2_smul_37056_comb, p2_sub_37057_comb);
  assign p2_sub_37155_comb = p2_sign_ext_36965_comb[47:32] - p2_sign_ext_36804_comb;
  assign p2_add_37201_comb = p1_sign_ext_36559 + {29'h0000_0000, {3{p1_sign_ext_36559[31]}}};
  assign p2_add_37206_comb = p1_sign_ext_36560 + {29'h0000_0000, {3{p1_sign_ext_36560[31]}}};
  assign p2_add_37211_comb = p1_sign_ext_36561 + {29'h0000_0000, {3{p1_sign_ext_36561[31]}}};
  assign p2_add_37216_comb = p1_sign_ext_36562 + {29'h0000_0000, {3{p1_sign_ext_36562[31]}}};
  assign p2_add_37221_comb = p1_sign_ext_36563 + {29'h0000_0000, {3{p1_sign_ext_36563[31]}}};
  assign p2_add_37226_comb = p1_sign_ext_36564 + {29'h0000_0000, {3{p1_sign_ext_36564[31]}}};
  assign p2_add_37231_comb = p1_sign_ext_36565 + {29'h0000_0000, {3{p1_sign_ext_36565[31]}}};
  assign p2_add_37236_comb = p1_sign_ext_36566 + {29'h0000_0000, {3{p1_sign_ext_36566[31]}}};
  assign p2_add_37240_comb = p2_sign_ext_36615_comb + {29'h0000_0000, {3{p2_sign_ext_36615_comb[31]}}};
  assign p2_add_37243_comb = p2_sign_ext_36616_comb + {29'h0000_0000, {3{p2_sign_ext_36616_comb[31]}}};
  assign p2_add_37246_comb = p2_sign_ext_36617_comb + {29'h0000_0000, {3{p2_sign_ext_36617_comb[31]}}};
  assign p2_add_37249_comb = p2_sign_ext_36618_comb + {29'h0000_0000, {3{p2_sign_ext_36618_comb[31]}}};
  assign p2_add_37252_comb = p2_sign_ext_36619_comb + {29'h0000_0000, {3{p2_sign_ext_36619_comb[31]}}};
  assign p2_add_37255_comb = p2_sign_ext_36620_comb + {29'h0000_0000, {3{p2_sign_ext_36620_comb[31]}}};
  assign p2_add_37258_comb = p2_sign_ext_36621_comb + {29'h0000_0000, {3{p2_sign_ext_36621_comb[31]}}};
  assign p2_add_37261_comb = p2_sign_ext_36622_comb + {29'h0000_0000, {3{p2_sign_ext_36622_comb[31]}}};
  assign p2_smul_37265_comb = smul47b_16b_x_31b(p1_neg_36543, 31'h2e8b_a2e9);
  assign p2_smul_37268_comb = smul47b_16b_x_31b(p1_neg_36544, 31'h2e8b_a2e9);
  assign p2_smul_37271_comb = smul47b_16b_x_31b(p1_neg_36545, 31'h2e8b_a2e9);
  assign p2_smul_37274_comb = smul47b_16b_x_31b(p1_neg_36546, 31'h2e8b_a2e9);
  assign p2_smul_37277_comb = smul47b_16b_x_31b(p1_neg_36547, 31'h2e8b_a2e9);
  assign p2_smul_37280_comb = smul47b_16b_x_31b(p1_neg_36548, 31'h2e8b_a2e9);
  assign p2_smul_37283_comb = smul47b_16b_x_31b(p1_neg_36549, 31'h2e8b_a2e9);
  assign p2_smul_37286_comb = smul47b_16b_x_31b(p1_neg_36550, 31'h2e8b_a2e9);
  assign p2_add_37471_comb = p1_sign_ext_36559 + {28'h000_0000, {4{p1_sign_ext_36559[31]}}};
  assign p2_add_37472_comb = p1_sign_ext_36560 + {28'h000_0000, {4{p1_sign_ext_36560[31]}}};
  assign p2_add_37473_comb = p1_sign_ext_36561 + {28'h000_0000, {4{p1_sign_ext_36561[31]}}};
  assign p2_add_37474_comb = p1_sign_ext_36562 + {28'h000_0000, {4{p1_sign_ext_36562[31]}}};
  assign p2_add_37475_comb = p1_sign_ext_36563 + {28'h000_0000, {4{p1_sign_ext_36563[31]}}};
  assign p2_add_37476_comb = p1_sign_ext_36564 + {28'h000_0000, {4{p1_sign_ext_36564[31]}}};
  assign p2_add_37477_comb = p1_sign_ext_36565 + {28'h000_0000, {4{p1_sign_ext_36565[31]}}};
  assign p2_add_37478_comb = p1_sign_ext_36566 + {28'h000_0000, {4{p1_sign_ext_36566[31]}}};
  assign p2_add_37479_comb = p2_sign_ext_36615_comb + {28'h000_0000, {4{p2_sign_ext_36615_comb[31]}}};
  assign p2_add_37480_comb = p2_sign_ext_36616_comb + {28'h000_0000, {4{p2_sign_ext_36616_comb[31]}}};
  assign p2_add_37481_comb = p2_sign_ext_36617_comb + {28'h000_0000, {4{p2_sign_ext_36617_comb[31]}}};
  assign p2_add_37482_comb = p2_sign_ext_36618_comb + {28'h000_0000, {4{p2_sign_ext_36618_comb[31]}}};
  assign p2_add_37483_comb = p2_sign_ext_36619_comb + {28'h000_0000, {4{p2_sign_ext_36619_comb[31]}}};
  assign p2_add_37484_comb = p2_sign_ext_36620_comb + {28'h000_0000, {4{p2_sign_ext_36620_comb[31]}}};
  assign p2_add_37485_comb = p2_sign_ext_36621_comb + {28'h000_0000, {4{p2_sign_ext_36621_comb[31]}}};
  assign p2_add_37486_comb = p2_sign_ext_36622_comb + {28'h000_0000, {4{p2_sign_ext_36622_comb[31]}}};
  assign p2_add_37535_comb = p1_neg_36543 + p2_smul_36847_comb;
  assign p2_add_37536_comb = p2_smul_36927_comb + p2_smul_37007_comb;
  assign p2_add_37537_comb = p1_neg_36544 + p2_smul_36852_comb;
  assign p2_add_37538_comb = p2_smul_36932_comb + p2_smul_37014_comb;
  assign p2_add_37539_comb = p1_neg_36545 + p2_smul_36857_comb;
  assign p2_add_37540_comb = p2_smul_36937_comb + p2_smul_37021_comb;
  assign p2_add_37541_comb = p1_neg_36546 + p2_smul_36862_comb;
  assign p2_add_37542_comb = p2_smul_36942_comb + p2_smul_37028_comb;
  assign p2_add_37543_comb = p1_neg_36547 + p2_smul_36867_comb;
  assign p2_add_37544_comb = p2_smul_36947_comb + p2_smul_37035_comb;
  assign p2_add_37545_comb = p1_neg_36548 + p2_smul_36872_comb;
  assign p2_add_37546_comb = p2_smul_36952_comb + p2_smul_37042_comb;
  assign p2_add_37547_comb = p1_neg_36549 + p2_smul_36877_comb;
  assign p2_add_37548_comb = p2_smul_36957_comb + p2_smul_37049_comb;
  assign p2_add_37549_comb = p1_neg_36550 + p2_smul_36882_comb;
  assign p2_add_37550_comb = p2_smul_36962_comb + p2_smul_37056_comb;
  assign p2_smul_37159_comb = smul16b_16b_x_16b(p2_smul_37063_comb, p2_sub_37064_comb);
  assign p2_sub_37160_comb = p2_sign_ext_36970_comb[47:32] - p2_sign_ext_36809_comb;
  assign p2_smul_37164_comb = smul16b_16b_x_16b(p2_smul_37070_comb, p2_sub_37071_comb);
  assign p2_sub_37165_comb = p2_sign_ext_36975_comb[47:32] - p2_sign_ext_36814_comb;
  assign p2_smul_37169_comb = smul16b_16b_x_16b(p2_smul_37077_comb, p2_sub_37078_comb);
  assign p2_sub_37170_comb = p2_sign_ext_36980_comb[47:32] - p2_sign_ext_36819_comb;
  assign p2_smul_37174_comb = smul16b_16b_x_16b(p2_smul_37084_comb, p2_sub_37085_comb);
  assign p2_sub_37175_comb = p2_sign_ext_36985_comb[47:32] - p2_sign_ext_36824_comb;
  assign p2_smul_37179_comb = smul16b_16b_x_16b(p2_smul_37091_comb, p2_sub_37092_comb);
  assign p2_sub_37180_comb = p2_sign_ext_36990_comb[47:32] - p2_sign_ext_36829_comb;
  assign p2_smul_37184_comb = smul16b_16b_x_16b(p2_smul_37098_comb, p2_sub_37099_comb);
  assign p2_sub_37185_comb = p2_sign_ext_36995_comb[47:32] - p2_sign_ext_36834_comb;
  assign p2_smul_37189_comb = smul16b_16b_x_16b(p2_smul_37105_comb, p2_sub_37106_comb);
  assign p2_sub_37190_comb = p2_sign_ext_37000_comb[47:32] - p2_sign_ext_36839_comb;
  assign p2_smul_37194_comb = smul16b_16b_x_16b(p2_smul_37112_comb, p2_sub_37113_comb);
  assign p2_sub_37195_comb = p2_sign_ext_37005_comb[47:32] - p2_sign_ext_36844_comb;
  assign p2_smul_37199_comb = smul16b_16b_x_16b(p2_smul_37119_comb, p2_sub_37120_comb);
  assign p2_sub_37200_comb = p2_sign_ext_37010_comb[49:34] - p2_sign_ext_36769_comb;
  assign p2_smul_37204_comb = smul16b_16b_x_16b(p2_smul_37124_comb, p2_sub_37125_comb);
  assign p2_sub_37205_comb = p2_sign_ext_37017_comb[49:34] - p2_sign_ext_36774_comb;
  assign p2_smul_37209_comb = smul16b_16b_x_16b(p2_smul_37129_comb, p2_sub_37130_comb);
  assign p2_sub_37210_comb = p2_sign_ext_37024_comb[49:34] - p2_sign_ext_36779_comb;
  assign p2_smul_37214_comb = smul16b_16b_x_16b(p2_smul_37134_comb, p2_sub_37135_comb);
  assign p2_sub_37215_comb = p2_sign_ext_37031_comb[49:34] - p2_sign_ext_36784_comb;
  assign p2_smul_37219_comb = smul16b_16b_x_16b(p2_smul_37139_comb, p2_sub_37140_comb);
  assign p2_sub_37220_comb = p2_sign_ext_37038_comb[49:34] - p2_sign_ext_36789_comb;
  assign p2_smul_37224_comb = smul16b_16b_x_16b(p2_smul_37144_comb, p2_sub_37145_comb);
  assign p2_sub_37225_comb = p2_sign_ext_37045_comb[49:34] - p2_sign_ext_36794_comb;
  assign p2_smul_37229_comb = smul16b_16b_x_16b(p2_smul_37149_comb, p2_sub_37150_comb);
  assign p2_sub_37230_comb = p2_sign_ext_37052_comb[49:34] - p2_sign_ext_36799_comb;
  assign p2_smul_37234_comb = smul16b_16b_x_16b(p2_smul_37154_comb, p2_sub_37155_comb);
  assign p2_sub_37235_comb = p2_sign_ext_37059_comb[49:34] - p2_sign_ext_36804_comb;
  assign p2_sub_37239_comb = p2_sign_ext_37066_comb[49:34] - p2_sign_ext_36809_comb;
  assign p2_sub_37242_comb = p2_sign_ext_37073_comb[49:34] - p2_sign_ext_36814_comb;
  assign p2_sub_37245_comb = p2_sign_ext_37080_comb[49:34] - p2_sign_ext_36819_comb;
  assign p2_sub_37248_comb = p2_sign_ext_37087_comb[49:34] - p2_sign_ext_36824_comb;
  assign p2_sub_37251_comb = p2_sign_ext_37094_comb[49:34] - p2_sign_ext_36829_comb;
  assign p2_sub_37254_comb = p2_sign_ext_37101_comb[49:34] - p2_sign_ext_36834_comb;
  assign p2_sub_37257_comb = p2_sign_ext_37108_comb[49:34] - p2_sign_ext_36839_comb;
  assign p2_sub_37260_comb = p2_sign_ext_37115_comb[49:34] - p2_sign_ext_36844_comb;
  assign p2_bit_slice_37263_comb = p2_add_37201_comb[18:3];
  assign p2_bit_slice_37266_comb = p2_add_37206_comb[18:3];
  assign p2_bit_slice_37269_comb = p2_add_37211_comb[18:3];
  assign p2_bit_slice_37272_comb = p2_add_37216_comb[18:3];
  assign p2_bit_slice_37275_comb = p2_add_37221_comb[18:3];
  assign p2_bit_slice_37278_comb = p2_add_37226_comb[18:3];
  assign p2_bit_slice_37281_comb = p2_add_37231_comb[18:3];
  assign p2_bit_slice_37284_comb = p2_add_37236_comb[18:3];
  assign p2_bit_slice_37287_comb = p2_add_37240_comb[18:3];
  assign p2_bit_slice_37289_comb = p2_add_37243_comb[18:3];
  assign p2_bit_slice_37291_comb = p2_add_37246_comb[18:3];
  assign p2_bit_slice_37293_comb = p2_add_37249_comb[18:3];
  assign p2_bit_slice_37295_comb = p2_add_37252_comb[18:3];
  assign p2_bit_slice_37297_comb = p2_add_37255_comb[18:3];
  assign p2_bit_slice_37299_comb = p2_add_37258_comb[18:3];
  assign p2_bit_slice_37301_comb = p2_add_37261_comb[18:3];
  assign p2_sub_37303_comb = p2_sign_ext_37202_comb[48:33] - p2_sign_ext_36769_comb;
  assign p2_bit_slice_37305_comb = p2_smul_37265_comb[46:33];
  assign p2_sub_37306_comb = p2_sign_ext_37207_comb[48:33] - p2_sign_ext_36774_comb;
  assign p2_bit_slice_37308_comb = p2_smul_37268_comb[46:33];
  assign p2_sub_37309_comb = p2_sign_ext_37212_comb[48:33] - p2_sign_ext_36779_comb;
  assign p2_bit_slice_37311_comb = p2_smul_37271_comb[46:33];
  assign p2_sub_37312_comb = p2_sign_ext_37217_comb[48:33] - p2_sign_ext_36784_comb;
  assign p2_bit_slice_37314_comb = p2_smul_37274_comb[46:33];
  assign p2_sub_37315_comb = p2_sign_ext_37222_comb[48:33] - p2_sign_ext_36789_comb;
  assign p2_bit_slice_37317_comb = p2_smul_37277_comb[46:33];
  assign p2_sub_37318_comb = p2_sign_ext_37227_comb[48:33] - p2_sign_ext_36794_comb;
  assign p2_bit_slice_37320_comb = p2_smul_37280_comb[46:33];
  assign p2_sub_37321_comb = p2_sign_ext_37232_comb[48:33] - p2_sign_ext_36799_comb;
  assign p2_bit_slice_37323_comb = p2_smul_37283_comb[46:33];
  assign p2_sub_37324_comb = p2_sign_ext_37237_comb[48:33] - p2_sign_ext_36804_comb;
  assign p2_bit_slice_37326_comb = p2_smul_37286_comb[46:33];
  assign p2_sub_37327_comb = p2_sign_ext_37241_comb[48:33] - p2_sign_ext_36809_comb;
  assign p2_sub_37329_comb = p2_sign_ext_37244_comb[48:33] - p2_sign_ext_36814_comb;
  assign p2_sub_37331_comb = p2_sign_ext_37247_comb[48:33] - p2_sign_ext_36819_comb;
  assign p2_sub_37333_comb = p2_sign_ext_37250_comb[48:33] - p2_sign_ext_36824_comb;
  assign p2_sub_37335_comb = p2_sign_ext_37253_comb[48:33] - p2_sign_ext_36829_comb;
  assign p2_sub_37337_comb = p2_sign_ext_37256_comb[48:33] - p2_sign_ext_36834_comb;
  assign p2_sub_37339_comb = p2_sign_ext_37259_comb[48:33] - p2_sign_ext_36839_comb;
  assign p2_sub_37341_comb = p2_sign_ext_37262_comb[48:33] - p2_sign_ext_36844_comb;
  assign p2_sub_37343_comb = p2_sign_ext_36850_comb[49:34] - p2_sign_ext_36769_comb;
  assign p2_sub_37344_comb = p2_sign_ext_36855_comb[49:34] - p2_sign_ext_36774_comb;
  assign p2_sub_37345_comb = p2_sign_ext_36860_comb[49:34] - p2_sign_ext_36779_comb;
  assign p2_sub_37346_comb = p2_sign_ext_36865_comb[49:34] - p2_sign_ext_36784_comb;
  assign p2_sub_37347_comb = p2_sign_ext_36870_comb[49:34] - p2_sign_ext_36789_comb;
  assign p2_sub_37348_comb = p2_sign_ext_36875_comb[49:34] - p2_sign_ext_36794_comb;
  assign p2_sub_37349_comb = p2_sign_ext_36880_comb[49:34] - p2_sign_ext_36799_comb;
  assign p2_sub_37350_comb = p2_sign_ext_36885_comb[49:34] - p2_sign_ext_36804_comb;
  assign p2_sub_37351_comb = p2_sign_ext_36890_comb[49:34] - p2_sign_ext_36809_comb;
  assign p2_sub_37352_comb = p2_sign_ext_36895_comb[49:34] - p2_sign_ext_36814_comb;
  assign p2_sub_37353_comb = p2_sign_ext_36900_comb[49:34] - p2_sign_ext_36819_comb;
  assign p2_sub_37354_comb = p2_sign_ext_36905_comb[49:34] - p2_sign_ext_36824_comb;
  assign p2_sub_37355_comb = p2_sign_ext_36910_comb[49:34] - p2_sign_ext_36829_comb;
  assign p2_sub_37356_comb = p2_sign_ext_36915_comb[49:34] - p2_sign_ext_36834_comb;
  assign p2_sub_37357_comb = p2_sign_ext_36920_comb[49:34] - p2_sign_ext_36839_comb;
  assign p2_sub_37358_comb = p2_sign_ext_36925_comb[49:34] - p2_sign_ext_36844_comb;
  assign p2_sub_37375_comb = p2_sign_ext_36930_comb[48:33] - p2_sign_ext_36769_comb;
  assign p2_sub_37376_comb = p2_sign_ext_36935_comb[48:33] - p2_sign_ext_36774_comb;
  assign p2_sub_37377_comb = p2_sign_ext_36940_comb[48:33] - p2_sign_ext_36779_comb;
  assign p2_sub_37378_comb = p2_sign_ext_36945_comb[48:33] - p2_sign_ext_36784_comb;
  assign p2_sub_37379_comb = p2_sign_ext_36950_comb[48:33] - p2_sign_ext_36789_comb;
  assign p2_sub_37380_comb = p2_sign_ext_36955_comb[48:33] - p2_sign_ext_36794_comb;
  assign p2_sub_37381_comb = p2_sign_ext_36960_comb[48:33] - p2_sign_ext_36799_comb;
  assign p2_sub_37382_comb = p2_sign_ext_36965_comb[48:33] - p2_sign_ext_36804_comb;
  assign p2_sub_37383_comb = p2_sign_ext_36970_comb[48:33] - p2_sign_ext_36809_comb;
  assign p2_sub_37384_comb = p2_sign_ext_36975_comb[48:33] - p2_sign_ext_36814_comb;
  assign p2_sub_37385_comb = p2_sign_ext_36980_comb[48:33] - p2_sign_ext_36819_comb;
  assign p2_sub_37386_comb = p2_sign_ext_36985_comb[48:33] - p2_sign_ext_36824_comb;
  assign p2_sub_37387_comb = p2_sign_ext_36990_comb[48:33] - p2_sign_ext_36829_comb;
  assign p2_sub_37388_comb = p2_sign_ext_36995_comb[48:33] - p2_sign_ext_36834_comb;
  assign p2_sub_37389_comb = p2_sign_ext_37000_comb[48:33] - p2_sign_ext_36839_comb;
  assign p2_sub_37390_comb = p2_sign_ext_37005_comb[48:33] - p2_sign_ext_36844_comb;
  assign p2_sub_37439_comb = p2_sign_ext_37010_comb[50:35] - p2_sign_ext_36769_comb;
  assign p2_sub_37441_comb = p2_sign_ext_37017_comb[50:35] - p2_sign_ext_36774_comb;
  assign p2_sub_37443_comb = p2_sign_ext_37024_comb[50:35] - p2_sign_ext_36779_comb;
  assign p2_sub_37445_comb = p2_sign_ext_37031_comb[50:35] - p2_sign_ext_36784_comb;
  assign p2_sub_37447_comb = p2_sign_ext_37038_comb[50:35] - p2_sign_ext_36789_comb;
  assign p2_sub_37449_comb = p2_sign_ext_37045_comb[50:35] - p2_sign_ext_36794_comb;
  assign p2_sub_37451_comb = p2_sign_ext_37052_comb[50:35] - p2_sign_ext_36799_comb;
  assign p2_sub_37453_comb = p2_sign_ext_37059_comb[50:35] - p2_sign_ext_36804_comb;
  assign p2_sub_37455_comb = p2_sign_ext_37066_comb[50:35] - p2_sign_ext_36809_comb;
  assign p2_sub_37457_comb = p2_sign_ext_37073_comb[50:35] - p2_sign_ext_36814_comb;
  assign p2_sub_37459_comb = p2_sign_ext_37080_comb[50:35] - p2_sign_ext_36819_comb;
  assign p2_sub_37461_comb = p2_sign_ext_37087_comb[50:35] - p2_sign_ext_36824_comb;
  assign p2_sub_37463_comb = p2_sign_ext_37094_comb[50:35] - p2_sign_ext_36829_comb;
  assign p2_sub_37465_comb = p2_sign_ext_37101_comb[50:35] - p2_sign_ext_36834_comb;
  assign p2_sub_37467_comb = p2_sign_ext_37108_comb[50:35] - p2_sign_ext_36839_comb;
  assign p2_sub_37469_comb = p2_sign_ext_37115_comb[50:35] - p2_sign_ext_36844_comb;
  assign p2_bit_slice_37487_comb = p2_add_37471_comb[19:4];
  assign p2_bit_slice_37488_comb = p2_add_37472_comb[19:4];
  assign p2_bit_slice_37489_comb = p2_add_37473_comb[19:4];
  assign p2_bit_slice_37490_comb = p2_add_37474_comb[19:4];
  assign p2_bit_slice_37491_comb = p2_add_37475_comb[19:4];
  assign p2_bit_slice_37492_comb = p2_add_37476_comb[19:4];
  assign p2_bit_slice_37493_comb = p2_add_37477_comb[19:4];
  assign p2_bit_slice_37494_comb = p2_add_37478_comb[19:4];
  assign p2_bit_slice_37495_comb = p2_add_37479_comb[19:4];
  assign p2_bit_slice_37496_comb = p2_add_37480_comb[19:4];
  assign p2_bit_slice_37497_comb = p2_add_37481_comb[19:4];
  assign p2_bit_slice_37498_comb = p2_add_37482_comb[19:4];
  assign p2_bit_slice_37499_comb = p2_add_37483_comb[19:4];
  assign p2_bit_slice_37500_comb = p2_add_37484_comb[19:4];
  assign p2_bit_slice_37501_comb = p2_add_37485_comb[19:4];
  assign p2_bit_slice_37502_comb = p2_add_37486_comb[19:4];
  assign p2_sub_37519_comb = p2_sign_ext_37202_comb[49:34] - p2_sign_ext_36769_comb;
  assign p2_sub_37520_comb = p2_sign_ext_37207_comb[49:34] - p2_sign_ext_36774_comb;
  assign p2_sub_37521_comb = p2_sign_ext_37212_comb[49:34] - p2_sign_ext_36779_comb;
  assign p2_sub_37522_comb = p2_sign_ext_37217_comb[49:34] - p2_sign_ext_36784_comb;
  assign p2_sub_37523_comb = p2_sign_ext_37222_comb[49:34] - p2_sign_ext_36789_comb;
  assign p2_sub_37524_comb = p2_sign_ext_37227_comb[49:34] - p2_sign_ext_36794_comb;
  assign p2_sub_37525_comb = p2_sign_ext_37232_comb[49:34] - p2_sign_ext_36799_comb;
  assign p2_sub_37526_comb = p2_sign_ext_37237_comb[49:34] - p2_sign_ext_36804_comb;
  assign p2_sub_37527_comb = p2_sign_ext_37241_comb[49:34] - p2_sign_ext_36809_comb;
  assign p2_sub_37528_comb = p2_sign_ext_37244_comb[49:34] - p2_sign_ext_36814_comb;
  assign p2_sub_37529_comb = p2_sign_ext_37247_comb[49:34] - p2_sign_ext_36819_comb;
  assign p2_sub_37530_comb = p2_sign_ext_37250_comb[49:34] - p2_sign_ext_36824_comb;
  assign p2_sub_37531_comb = p2_sign_ext_37253_comb[49:34] - p2_sign_ext_36829_comb;
  assign p2_sub_37532_comb = p2_sign_ext_37256_comb[49:34] - p2_sign_ext_36834_comb;
  assign p2_sub_37533_comb = p2_sign_ext_37259_comb[49:34] - p2_sign_ext_36839_comb;
  assign p2_sub_37534_comb = p2_sign_ext_37262_comb[49:34] - p2_sign_ext_36844_comb;
  assign p2_add_37551_comb = p1_neg_36551 + p2_smul_36887_comb;
  assign p2_add_37552_comb = p2_smul_36967_comb + p2_smul_37063_comb;
  assign p2_add_37553_comb = p1_neg_36552 + p2_smul_36892_comb;
  assign p2_add_37554_comb = p2_smul_36972_comb + p2_smul_37070_comb;
  assign p2_add_37555_comb = p1_neg_36553 + p2_smul_36897_comb;
  assign p2_add_37556_comb = p2_smul_36977_comb + p2_smul_37077_comb;
  assign p2_add_37557_comb = p1_neg_36554 + p2_smul_36902_comb;
  assign p2_add_37558_comb = p2_smul_36982_comb + p2_smul_37084_comb;
  assign p2_add_37559_comb = p1_neg_36555 + p2_smul_36907_comb;
  assign p2_add_37560_comb = p2_smul_36987_comb + p2_smul_37091_comb;
  assign p2_add_37561_comb = p1_neg_36556 + p2_smul_36912_comb;
  assign p2_add_37562_comb = p2_smul_36992_comb + p2_smul_37098_comb;
  assign p2_add_37563_comb = p1_neg_36557 + p2_smul_36917_comb;
  assign p2_add_37564_comb = p2_smul_36997_comb + p2_smul_37105_comb;
  assign p2_add_37565_comb = p1_neg_36558 + p2_smul_36922_comb;
  assign p2_add_37566_comb = p2_smul_37002_comb + p2_smul_37112_comb;
  assign p2_add_37567_comb = p2_add_37535_comb + p2_add_37536_comb;
  assign p2_add_37568_comb = p2_add_37537_comb + p2_add_37538_comb;
  assign p2_add_37569_comb = p2_add_37539_comb + p2_add_37540_comb;
  assign p2_add_37570_comb = p2_add_37541_comb + p2_add_37542_comb;
  assign p2_add_37571_comb = p2_add_37543_comb + p2_add_37544_comb;
  assign p2_add_37572_comb = p2_add_37545_comb + p2_add_37546_comb;
  assign p2_add_37573_comb = p2_add_37547_comb + p2_add_37548_comb;
  assign p2_add_37574_comb = p2_add_37549_comb + p2_add_37550_comb;

  // Registers for pipe stage 2:
  reg [15:0] p2_neg_36543;
  reg [15:0] p2_neg_36544;
  reg [15:0] p2_neg_36545;
  reg [15:0] p2_neg_36546;
  reg [15:0] p2_neg_36547;
  reg [15:0] p2_neg_36548;
  reg [15:0] p2_neg_36549;
  reg [15:0] p2_neg_36550;
  reg [15:0] p2_neg_36551;
  reg [15:0] p2_neg_36552;
  reg [15:0] p2_neg_36553;
  reg [15:0] p2_neg_36554;
  reg [15:0] p2_neg_36555;
  reg [15:0] p2_neg_36556;
  reg [15:0] p2_neg_36557;
  reg [15:0] p2_neg_36558;
  reg [15:0] p2_sign_ext_36769;
  reg [15:0] p2_sign_ext_36774;
  reg [15:0] p2_sign_ext_36779;
  reg [15:0] p2_sign_ext_36784;
  reg [15:0] p2_sign_ext_36789;
  reg [15:0] p2_sign_ext_36794;
  reg [15:0] p2_sign_ext_36799;
  reg [15:0] p2_sign_ext_36804;
  reg [15:0] p2_sign_ext_36809;
  reg [15:0] p2_sign_ext_36814;
  reg [15:0] p2_sign_ext_36819;
  reg [15:0] p2_sign_ext_36824;
  reg [15:0] p2_sign_ext_36829;
  reg [15:0] p2_sign_ext_36834;
  reg [15:0] p2_sign_ext_36839;
  reg [15:0] p2_sign_ext_36844;
  reg [15:0] p2_smul_37119;
  reg [15:0] p2_smul_37124;
  reg [15:0] p2_smul_37129;
  reg [15:0] p2_smul_37134;
  reg [15:0] p2_smul_37139;
  reg [15:0] p2_smul_37144;
  reg [15:0] p2_smul_37149;
  reg [15:0] p2_smul_37154;
  reg [15:0] p2_smul_37159;
  reg [15:0] p2_sub_37160;
  reg [15:0] p2_smul_37164;
  reg [15:0] p2_sub_37165;
  reg [15:0] p2_smul_37169;
  reg [15:0] p2_sub_37170;
  reg [15:0] p2_smul_37174;
  reg [15:0] p2_sub_37175;
  reg [15:0] p2_smul_37179;
  reg [15:0] p2_sub_37180;
  reg [15:0] p2_smul_37184;
  reg [15:0] p2_sub_37185;
  reg [15:0] p2_smul_37189;
  reg [15:0] p2_sub_37190;
  reg [15:0] p2_smul_37194;
  reg [15:0] p2_sub_37195;
  reg [15:0] p2_smul_37199;
  reg [15:0] p2_sub_37200;
  reg [15:0] p2_smul_37204;
  reg [15:0] p2_sub_37205;
  reg [15:0] p2_smul_37209;
  reg [15:0] p2_sub_37210;
  reg [15:0] p2_smul_37214;
  reg [15:0] p2_sub_37215;
  reg [15:0] p2_smul_37219;
  reg [15:0] p2_sub_37220;
  reg [15:0] p2_smul_37224;
  reg [15:0] p2_sub_37225;
  reg [15:0] p2_smul_37229;
  reg [15:0] p2_sub_37230;
  reg [15:0] p2_smul_37234;
  reg [15:0] p2_sub_37235;
  reg [15:0] p2_sub_37239;
  reg [15:0] p2_sub_37242;
  reg [15:0] p2_sub_37245;
  reg [15:0] p2_sub_37248;
  reg [15:0] p2_sub_37251;
  reg [15:0] p2_sub_37254;
  reg [15:0] p2_sub_37257;
  reg [15:0] p2_sub_37260;
  reg [15:0] p2_bit_slice_37263;
  reg [15:0] p2_bit_slice_37266;
  reg [15:0] p2_bit_slice_37269;
  reg [15:0] p2_bit_slice_37272;
  reg [15:0] p2_bit_slice_37275;
  reg [15:0] p2_bit_slice_37278;
  reg [15:0] p2_bit_slice_37281;
  reg [15:0] p2_bit_slice_37284;
  reg [15:0] p2_bit_slice_37287;
  reg [15:0] p2_bit_slice_37289;
  reg [15:0] p2_bit_slice_37291;
  reg [15:0] p2_bit_slice_37293;
  reg [15:0] p2_bit_slice_37295;
  reg [15:0] p2_bit_slice_37297;
  reg [15:0] p2_bit_slice_37299;
  reg [15:0] p2_bit_slice_37301;
  reg [15:0] p2_sub_37303;
  reg [13:0] p2_bit_slice_37305;
  reg [15:0] p2_sub_37306;
  reg [13:0] p2_bit_slice_37308;
  reg [15:0] p2_sub_37309;
  reg [13:0] p2_bit_slice_37311;
  reg [15:0] p2_sub_37312;
  reg [13:0] p2_bit_slice_37314;
  reg [15:0] p2_sub_37315;
  reg [13:0] p2_bit_slice_37317;
  reg [15:0] p2_sub_37318;
  reg [13:0] p2_bit_slice_37320;
  reg [15:0] p2_sub_37321;
  reg [13:0] p2_bit_slice_37323;
  reg [15:0] p2_sub_37324;
  reg [13:0] p2_bit_slice_37326;
  reg [15:0] p2_sub_37327;
  reg [15:0] p2_sub_37329;
  reg [15:0] p2_sub_37331;
  reg [15:0] p2_sub_37333;
  reg [15:0] p2_sub_37335;
  reg [15:0] p2_sub_37337;
  reg [15:0] p2_sub_37339;
  reg [15:0] p2_sub_37341;
  reg [15:0] p2_sub_37343;
  reg [15:0] p2_sub_37344;
  reg [15:0] p2_sub_37345;
  reg [15:0] p2_sub_37346;
  reg [15:0] p2_sub_37347;
  reg [15:0] p2_sub_37348;
  reg [15:0] p2_sub_37349;
  reg [15:0] p2_sub_37350;
  reg [15:0] p2_sub_37351;
  reg [15:0] p2_sub_37352;
  reg [15:0] p2_sub_37353;
  reg [15:0] p2_sub_37354;
  reg [15:0] p2_sub_37355;
  reg [15:0] p2_sub_37356;
  reg [15:0] p2_sub_37357;
  reg [15:0] p2_sub_37358;
  reg [15:0] p2_sub_37375;
  reg [15:0] p2_sub_37376;
  reg [15:0] p2_sub_37377;
  reg [15:0] p2_sub_37378;
  reg [15:0] p2_sub_37379;
  reg [15:0] p2_sub_37380;
  reg [15:0] p2_sub_37381;
  reg [15:0] p2_sub_37382;
  reg [15:0] p2_sub_37383;
  reg [15:0] p2_sub_37384;
  reg [15:0] p2_sub_37385;
  reg [15:0] p2_sub_37386;
  reg [15:0] p2_sub_37387;
  reg [15:0] p2_sub_37388;
  reg [15:0] p2_sub_37389;
  reg [15:0] p2_sub_37390;
  reg [15:0] p2_sub_37439;
  reg [15:0] p2_sub_37441;
  reg [15:0] p2_sub_37443;
  reg [15:0] p2_sub_37445;
  reg [15:0] p2_sub_37447;
  reg [15:0] p2_sub_37449;
  reg [15:0] p2_sub_37451;
  reg [15:0] p2_sub_37453;
  reg [15:0] p2_sub_37455;
  reg [15:0] p2_sub_37457;
  reg [15:0] p2_sub_37459;
  reg [15:0] p2_sub_37461;
  reg [15:0] p2_sub_37463;
  reg [15:0] p2_sub_37465;
  reg [15:0] p2_sub_37467;
  reg [15:0] p2_sub_37469;
  reg [15:0] p2_bit_slice_37487;
  reg [15:0] p2_bit_slice_37488;
  reg [15:0] p2_bit_slice_37489;
  reg [15:0] p2_bit_slice_37490;
  reg [15:0] p2_bit_slice_37491;
  reg [15:0] p2_bit_slice_37492;
  reg [15:0] p2_bit_slice_37493;
  reg [15:0] p2_bit_slice_37494;
  reg [15:0] p2_bit_slice_37495;
  reg [15:0] p2_bit_slice_37496;
  reg [15:0] p2_bit_slice_37497;
  reg [15:0] p2_bit_slice_37498;
  reg [15:0] p2_bit_slice_37499;
  reg [15:0] p2_bit_slice_37500;
  reg [15:0] p2_bit_slice_37501;
  reg [15:0] p2_bit_slice_37502;
  reg [15:0] p2_sub_37519;
  reg [15:0] p2_sub_37520;
  reg [15:0] p2_sub_37521;
  reg [15:0] p2_sub_37522;
  reg [15:0] p2_sub_37523;
  reg [15:0] p2_sub_37524;
  reg [15:0] p2_sub_37525;
  reg [15:0] p2_sub_37526;
  reg [15:0] p2_sub_37527;
  reg [15:0] p2_sub_37528;
  reg [15:0] p2_sub_37529;
  reg [15:0] p2_sub_37530;
  reg [15:0] p2_sub_37531;
  reg [15:0] p2_sub_37532;
  reg [15:0] p2_sub_37533;
  reg [15:0] p2_sub_37534;
  reg [15:0] p2_add_37551;
  reg [15:0] p2_add_37552;
  reg [15:0] p2_add_37553;
  reg [15:0] p2_add_37554;
  reg [15:0] p2_add_37555;
  reg [15:0] p2_add_37556;
  reg [15:0] p2_add_37557;
  reg [15:0] p2_add_37558;
  reg [15:0] p2_add_37559;
  reg [15:0] p2_add_37560;
  reg [15:0] p2_add_37561;
  reg [15:0] p2_add_37562;
  reg [15:0] p2_add_37563;
  reg [15:0] p2_add_37564;
  reg [15:0] p2_add_37565;
  reg [15:0] p2_add_37566;
  reg [15:0] p2_add_37567;
  reg [15:0] p2_add_37568;
  reg [15:0] p2_add_37569;
  reg [15:0] p2_add_37570;
  reg [15:0] p2_add_37571;
  reg [15:0] p2_add_37572;
  reg [15:0] p2_add_37573;
  reg [15:0] p2_add_37574;
  always_ff @ (posedge clk) begin
    p2_neg_36543 <= p1_neg_36543;
    p2_neg_36544 <= p1_neg_36544;
    p2_neg_36545 <= p1_neg_36545;
    p2_neg_36546 <= p1_neg_36546;
    p2_neg_36547 <= p1_neg_36547;
    p2_neg_36548 <= p1_neg_36548;
    p2_neg_36549 <= p1_neg_36549;
    p2_neg_36550 <= p1_neg_36550;
    p2_neg_36551 <= p1_neg_36551;
    p2_neg_36552 <= p1_neg_36552;
    p2_neg_36553 <= p1_neg_36553;
    p2_neg_36554 <= p1_neg_36554;
    p2_neg_36555 <= p1_neg_36555;
    p2_neg_36556 <= p1_neg_36556;
    p2_neg_36557 <= p1_neg_36557;
    p2_neg_36558 <= p1_neg_36558;
    p2_sign_ext_36769 <= p2_sign_ext_36769_comb;
    p2_sign_ext_36774 <= p2_sign_ext_36774_comb;
    p2_sign_ext_36779 <= p2_sign_ext_36779_comb;
    p2_sign_ext_36784 <= p2_sign_ext_36784_comb;
    p2_sign_ext_36789 <= p2_sign_ext_36789_comb;
    p2_sign_ext_36794 <= p2_sign_ext_36794_comb;
    p2_sign_ext_36799 <= p2_sign_ext_36799_comb;
    p2_sign_ext_36804 <= p2_sign_ext_36804_comb;
    p2_sign_ext_36809 <= p2_sign_ext_36809_comb;
    p2_sign_ext_36814 <= p2_sign_ext_36814_comb;
    p2_sign_ext_36819 <= p2_sign_ext_36819_comb;
    p2_sign_ext_36824 <= p2_sign_ext_36824_comb;
    p2_sign_ext_36829 <= p2_sign_ext_36829_comb;
    p2_sign_ext_36834 <= p2_sign_ext_36834_comb;
    p2_sign_ext_36839 <= p2_sign_ext_36839_comb;
    p2_sign_ext_36844 <= p2_sign_ext_36844_comb;
    p2_smul_37119 <= p2_smul_37119_comb;
    p2_smul_37124 <= p2_smul_37124_comb;
    p2_smul_37129 <= p2_smul_37129_comb;
    p2_smul_37134 <= p2_smul_37134_comb;
    p2_smul_37139 <= p2_smul_37139_comb;
    p2_smul_37144 <= p2_smul_37144_comb;
    p2_smul_37149 <= p2_smul_37149_comb;
    p2_smul_37154 <= p2_smul_37154_comb;
    p2_smul_37159 <= p2_smul_37159_comb;
    p2_sub_37160 <= p2_sub_37160_comb;
    p2_smul_37164 <= p2_smul_37164_comb;
    p2_sub_37165 <= p2_sub_37165_comb;
    p2_smul_37169 <= p2_smul_37169_comb;
    p2_sub_37170 <= p2_sub_37170_comb;
    p2_smul_37174 <= p2_smul_37174_comb;
    p2_sub_37175 <= p2_sub_37175_comb;
    p2_smul_37179 <= p2_smul_37179_comb;
    p2_sub_37180 <= p2_sub_37180_comb;
    p2_smul_37184 <= p2_smul_37184_comb;
    p2_sub_37185 <= p2_sub_37185_comb;
    p2_smul_37189 <= p2_smul_37189_comb;
    p2_sub_37190 <= p2_sub_37190_comb;
    p2_smul_37194 <= p2_smul_37194_comb;
    p2_sub_37195 <= p2_sub_37195_comb;
    p2_smul_37199 <= p2_smul_37199_comb;
    p2_sub_37200 <= p2_sub_37200_comb;
    p2_smul_37204 <= p2_smul_37204_comb;
    p2_sub_37205 <= p2_sub_37205_comb;
    p2_smul_37209 <= p2_smul_37209_comb;
    p2_sub_37210 <= p2_sub_37210_comb;
    p2_smul_37214 <= p2_smul_37214_comb;
    p2_sub_37215 <= p2_sub_37215_comb;
    p2_smul_37219 <= p2_smul_37219_comb;
    p2_sub_37220 <= p2_sub_37220_comb;
    p2_smul_37224 <= p2_smul_37224_comb;
    p2_sub_37225 <= p2_sub_37225_comb;
    p2_smul_37229 <= p2_smul_37229_comb;
    p2_sub_37230 <= p2_sub_37230_comb;
    p2_smul_37234 <= p2_smul_37234_comb;
    p2_sub_37235 <= p2_sub_37235_comb;
    p2_sub_37239 <= p2_sub_37239_comb;
    p2_sub_37242 <= p2_sub_37242_comb;
    p2_sub_37245 <= p2_sub_37245_comb;
    p2_sub_37248 <= p2_sub_37248_comb;
    p2_sub_37251 <= p2_sub_37251_comb;
    p2_sub_37254 <= p2_sub_37254_comb;
    p2_sub_37257 <= p2_sub_37257_comb;
    p2_sub_37260 <= p2_sub_37260_comb;
    p2_bit_slice_37263 <= p2_bit_slice_37263_comb;
    p2_bit_slice_37266 <= p2_bit_slice_37266_comb;
    p2_bit_slice_37269 <= p2_bit_slice_37269_comb;
    p2_bit_slice_37272 <= p2_bit_slice_37272_comb;
    p2_bit_slice_37275 <= p2_bit_slice_37275_comb;
    p2_bit_slice_37278 <= p2_bit_slice_37278_comb;
    p2_bit_slice_37281 <= p2_bit_slice_37281_comb;
    p2_bit_slice_37284 <= p2_bit_slice_37284_comb;
    p2_bit_slice_37287 <= p2_bit_slice_37287_comb;
    p2_bit_slice_37289 <= p2_bit_slice_37289_comb;
    p2_bit_slice_37291 <= p2_bit_slice_37291_comb;
    p2_bit_slice_37293 <= p2_bit_slice_37293_comb;
    p2_bit_slice_37295 <= p2_bit_slice_37295_comb;
    p2_bit_slice_37297 <= p2_bit_slice_37297_comb;
    p2_bit_slice_37299 <= p2_bit_slice_37299_comb;
    p2_bit_slice_37301 <= p2_bit_slice_37301_comb;
    p2_sub_37303 <= p2_sub_37303_comb;
    p2_bit_slice_37305 <= p2_bit_slice_37305_comb;
    p2_sub_37306 <= p2_sub_37306_comb;
    p2_bit_slice_37308 <= p2_bit_slice_37308_comb;
    p2_sub_37309 <= p2_sub_37309_comb;
    p2_bit_slice_37311 <= p2_bit_slice_37311_comb;
    p2_sub_37312 <= p2_sub_37312_comb;
    p2_bit_slice_37314 <= p2_bit_slice_37314_comb;
    p2_sub_37315 <= p2_sub_37315_comb;
    p2_bit_slice_37317 <= p2_bit_slice_37317_comb;
    p2_sub_37318 <= p2_sub_37318_comb;
    p2_bit_slice_37320 <= p2_bit_slice_37320_comb;
    p2_sub_37321 <= p2_sub_37321_comb;
    p2_bit_slice_37323 <= p2_bit_slice_37323_comb;
    p2_sub_37324 <= p2_sub_37324_comb;
    p2_bit_slice_37326 <= p2_bit_slice_37326_comb;
    p2_sub_37327 <= p2_sub_37327_comb;
    p2_sub_37329 <= p2_sub_37329_comb;
    p2_sub_37331 <= p2_sub_37331_comb;
    p2_sub_37333 <= p2_sub_37333_comb;
    p2_sub_37335 <= p2_sub_37335_comb;
    p2_sub_37337 <= p2_sub_37337_comb;
    p2_sub_37339 <= p2_sub_37339_comb;
    p2_sub_37341 <= p2_sub_37341_comb;
    p2_sub_37343 <= p2_sub_37343_comb;
    p2_sub_37344 <= p2_sub_37344_comb;
    p2_sub_37345 <= p2_sub_37345_comb;
    p2_sub_37346 <= p2_sub_37346_comb;
    p2_sub_37347 <= p2_sub_37347_comb;
    p2_sub_37348 <= p2_sub_37348_comb;
    p2_sub_37349 <= p2_sub_37349_comb;
    p2_sub_37350 <= p2_sub_37350_comb;
    p2_sub_37351 <= p2_sub_37351_comb;
    p2_sub_37352 <= p2_sub_37352_comb;
    p2_sub_37353 <= p2_sub_37353_comb;
    p2_sub_37354 <= p2_sub_37354_comb;
    p2_sub_37355 <= p2_sub_37355_comb;
    p2_sub_37356 <= p2_sub_37356_comb;
    p2_sub_37357 <= p2_sub_37357_comb;
    p2_sub_37358 <= p2_sub_37358_comb;
    p2_sub_37375 <= p2_sub_37375_comb;
    p2_sub_37376 <= p2_sub_37376_comb;
    p2_sub_37377 <= p2_sub_37377_comb;
    p2_sub_37378 <= p2_sub_37378_comb;
    p2_sub_37379 <= p2_sub_37379_comb;
    p2_sub_37380 <= p2_sub_37380_comb;
    p2_sub_37381 <= p2_sub_37381_comb;
    p2_sub_37382 <= p2_sub_37382_comb;
    p2_sub_37383 <= p2_sub_37383_comb;
    p2_sub_37384 <= p2_sub_37384_comb;
    p2_sub_37385 <= p2_sub_37385_comb;
    p2_sub_37386 <= p2_sub_37386_comb;
    p2_sub_37387 <= p2_sub_37387_comb;
    p2_sub_37388 <= p2_sub_37388_comb;
    p2_sub_37389 <= p2_sub_37389_comb;
    p2_sub_37390 <= p2_sub_37390_comb;
    p2_sub_37439 <= p2_sub_37439_comb;
    p2_sub_37441 <= p2_sub_37441_comb;
    p2_sub_37443 <= p2_sub_37443_comb;
    p2_sub_37445 <= p2_sub_37445_comb;
    p2_sub_37447 <= p2_sub_37447_comb;
    p2_sub_37449 <= p2_sub_37449_comb;
    p2_sub_37451 <= p2_sub_37451_comb;
    p2_sub_37453 <= p2_sub_37453_comb;
    p2_sub_37455 <= p2_sub_37455_comb;
    p2_sub_37457 <= p2_sub_37457_comb;
    p2_sub_37459 <= p2_sub_37459_comb;
    p2_sub_37461 <= p2_sub_37461_comb;
    p2_sub_37463 <= p2_sub_37463_comb;
    p2_sub_37465 <= p2_sub_37465_comb;
    p2_sub_37467 <= p2_sub_37467_comb;
    p2_sub_37469 <= p2_sub_37469_comb;
    p2_bit_slice_37487 <= p2_bit_slice_37487_comb;
    p2_bit_slice_37488 <= p2_bit_slice_37488_comb;
    p2_bit_slice_37489 <= p2_bit_slice_37489_comb;
    p2_bit_slice_37490 <= p2_bit_slice_37490_comb;
    p2_bit_slice_37491 <= p2_bit_slice_37491_comb;
    p2_bit_slice_37492 <= p2_bit_slice_37492_comb;
    p2_bit_slice_37493 <= p2_bit_slice_37493_comb;
    p2_bit_slice_37494 <= p2_bit_slice_37494_comb;
    p2_bit_slice_37495 <= p2_bit_slice_37495_comb;
    p2_bit_slice_37496 <= p2_bit_slice_37496_comb;
    p2_bit_slice_37497 <= p2_bit_slice_37497_comb;
    p2_bit_slice_37498 <= p2_bit_slice_37498_comb;
    p2_bit_slice_37499 <= p2_bit_slice_37499_comb;
    p2_bit_slice_37500 <= p2_bit_slice_37500_comb;
    p2_bit_slice_37501 <= p2_bit_slice_37501_comb;
    p2_bit_slice_37502 <= p2_bit_slice_37502_comb;
    p2_sub_37519 <= p2_sub_37519_comb;
    p2_sub_37520 <= p2_sub_37520_comb;
    p2_sub_37521 <= p2_sub_37521_comb;
    p2_sub_37522 <= p2_sub_37522_comb;
    p2_sub_37523 <= p2_sub_37523_comb;
    p2_sub_37524 <= p2_sub_37524_comb;
    p2_sub_37525 <= p2_sub_37525_comb;
    p2_sub_37526 <= p2_sub_37526_comb;
    p2_sub_37527 <= p2_sub_37527_comb;
    p2_sub_37528 <= p2_sub_37528_comb;
    p2_sub_37529 <= p2_sub_37529_comb;
    p2_sub_37530 <= p2_sub_37530_comb;
    p2_sub_37531 <= p2_sub_37531_comb;
    p2_sub_37532 <= p2_sub_37532_comb;
    p2_sub_37533 <= p2_sub_37533_comb;
    p2_sub_37534 <= p2_sub_37534_comb;
    p2_add_37551 <= p2_add_37551_comb;
    p2_add_37552 <= p2_add_37552_comb;
    p2_add_37553 <= p2_add_37553_comb;
    p2_add_37554 <= p2_add_37554_comb;
    p2_add_37555 <= p2_add_37555_comb;
    p2_add_37556 <= p2_add_37556_comb;
    p2_add_37557 <= p2_add_37557_comb;
    p2_add_37558 <= p2_add_37558_comb;
    p2_add_37559 <= p2_add_37559_comb;
    p2_add_37560 <= p2_add_37560_comb;
    p2_add_37561 <= p2_add_37561_comb;
    p2_add_37562 <= p2_add_37562_comb;
    p2_add_37563 <= p2_add_37563_comb;
    p2_add_37564 <= p2_add_37564_comb;
    p2_add_37565 <= p2_add_37565_comb;
    p2_add_37566 <= p2_add_37566_comb;
    p2_add_37567 <= p2_add_37567_comb;
    p2_add_37568 <= p2_add_37568_comb;
    p2_add_37569 <= p2_add_37569_comb;
    p2_add_37570 <= p2_add_37570_comb;
    p2_add_37571 <= p2_add_37571_comb;
    p2_add_37572 <= p2_add_37572_comb;
    p2_add_37573 <= p2_add_37573_comb;
    p2_add_37574 <= p2_add_37574_comb;
  end

  // ===== Pipe stage 3:
  wire [15:0] p3_smul_38023_comb;
  wire [15:0] p3_smul_38025_comb;
  wire [15:0] p3_smul_38027_comb;
  wire [15:0] p3_smul_38029_comb;
  wire [15:0] p3_smul_38031_comb;
  wire [15:0] p3_smul_38033_comb;
  wire [15:0] p3_smul_38035_comb;
  wire [15:0] p3_smul_38037_comb;
  wire [15:0] p3_smul_38039_comb;
  wire [15:0] p3_smul_38040_comb;
  wire [15:0] p3_smul_38041_comb;
  wire [15:0] p3_smul_38042_comb;
  wire [15:0] p3_smul_38043_comb;
  wire [15:0] p3_smul_38044_comb;
  wire [15:0] p3_smul_38045_comb;
  wire [15:0] p3_smul_38046_comb;
  wire [15:0] p3_smul_38047_comb;
  wire [46:0] p3_smul_38048_comb;
  wire [15:0] p3_smul_38049_comb;
  wire [46:0] p3_smul_38050_comb;
  wire [15:0] p3_smul_38051_comb;
  wire [46:0] p3_smul_38052_comb;
  wire [15:0] p3_smul_38053_comb;
  wire [46:0] p3_smul_38054_comb;
  wire [15:0] p3_smul_38055_comb;
  wire [46:0] p3_smul_38056_comb;
  wire [15:0] p3_smul_38057_comb;
  wire [46:0] p3_smul_38058_comb;
  wire [15:0] p3_smul_38059_comb;
  wire [46:0] p3_smul_38060_comb;
  wire [15:0] p3_smul_38061_comb;
  wire [46:0] p3_smul_38062_comb;
  wire [15:0] p3_smul_38063_comb;
  wire [15:0] p3_smul_38065_comb;
  wire [15:0] p3_smul_38067_comb;
  wire [15:0] p3_smul_38069_comb;
  wire [15:0] p3_smul_38071_comb;
  wire [15:0] p3_smul_38073_comb;
  wire [15:0] p3_smul_38075_comb;
  wire [15:0] p3_smul_38077_comb;
  wire [15:0] p3_smul_38079_comb;
  wire [13:0] p3_bit_slice_38080_comb;
  wire [15:0] p3_smul_38082_comb;
  wire [13:0] p3_bit_slice_38083_comb;
  wire [15:0] p3_smul_38085_comb;
  wire [13:0] p3_bit_slice_38086_comb;
  wire [15:0] p3_smul_38088_comb;
  wire [13:0] p3_bit_slice_38089_comb;
  wire [15:0] p3_smul_38091_comb;
  wire [13:0] p3_bit_slice_38092_comb;
  wire [15:0] p3_smul_38094_comb;
  wire [13:0] p3_bit_slice_38095_comb;
  wire [15:0] p3_smul_38097_comb;
  wire [13:0] p3_bit_slice_38098_comb;
  wire [15:0] p3_smul_38100_comb;
  wire [13:0] p3_bit_slice_38101_comb;
  wire [15:0] p3_smul_38103_comb;
  wire [47:0] p3_smul_38105_comb;
  wire [15:0] p3_smul_38106_comb;
  wire [47:0] p3_smul_38108_comb;
  wire [15:0] p3_smul_38109_comb;
  wire [47:0] p3_smul_38111_comb;
  wire [15:0] p3_smul_38112_comb;
  wire [47:0] p3_smul_38114_comb;
  wire [15:0] p3_smul_38115_comb;
  wire [47:0] p3_smul_38117_comb;
  wire [15:0] p3_smul_38118_comb;
  wire [47:0] p3_smul_38120_comb;
  wire [15:0] p3_smul_38121_comb;
  wire [47:0] p3_smul_38123_comb;
  wire [15:0] p3_smul_38124_comb;
  wire [47:0] p3_smul_38126_comb;
  wire [15:0] p3_smul_38127_comb;
  wire [47:0] p3_smul_38129_comb;
  wire [15:0] p3_smul_38130_comb;
  wire [47:0] p3_smul_38132_comb;
  wire [15:0] p3_smul_38133_comb;
  wire [47:0] p3_smul_38135_comb;
  wire [15:0] p3_smul_38136_comb;
  wire [47:0] p3_smul_38138_comb;
  wire [15:0] p3_smul_38139_comb;
  wire [47:0] p3_smul_38141_comb;
  wire [15:0] p3_smul_38142_comb;
  wire [47:0] p3_smul_38144_comb;
  wire [15:0] p3_smul_38145_comb;
  wire [47:0] p3_smul_38147_comb;
  wire [15:0] p3_smul_38148_comb;
  wire [47:0] p3_smul_38150_comb;
  wire [15:0] p3_smul_38151_comb;
  wire [15:0] p3_sub_38152_comb;
  wire [13:0] p3_bit_slice_38153_comb;
  wire [15:0] p3_smul_38155_comb;
  wire [15:0] p3_sub_38156_comb;
  wire [13:0] p3_bit_slice_38157_comb;
  wire [15:0] p3_smul_38159_comb;
  wire [15:0] p3_sub_38160_comb;
  wire [13:0] p3_bit_slice_38161_comb;
  wire [15:0] p3_smul_38163_comb;
  wire [15:0] p3_sub_38164_comb;
  wire [13:0] p3_bit_slice_38165_comb;
  wire [15:0] p3_smul_38167_comb;
  wire [15:0] p3_sub_38168_comb;
  wire [13:0] p3_bit_slice_38169_comb;
  wire [15:0] p3_smul_38171_comb;
  wire [15:0] p3_sub_38172_comb;
  wire [13:0] p3_bit_slice_38173_comb;
  wire [15:0] p3_smul_38175_comb;
  wire [15:0] p3_sub_38176_comb;
  wire [13:0] p3_bit_slice_38177_comb;
  wire [15:0] p3_smul_38179_comb;
  wire [15:0] p3_sub_38180_comb;
  wire [13:0] p3_bit_slice_38181_comb;
  wire [15:0] p3_smul_38183_comb;
  wire [15:0] p3_sub_38184_comb;
  wire [13:0] p3_bit_slice_38185_comb;
  wire [15:0] p3_smul_38187_comb;
  wire [15:0] p3_sub_38188_comb;
  wire [13:0] p3_bit_slice_38189_comb;
  wire [15:0] p3_smul_38191_comb;
  wire [15:0] p3_sub_38192_comb;
  wire [13:0] p3_bit_slice_38193_comb;
  wire [15:0] p3_smul_38195_comb;
  wire [15:0] p3_sub_38196_comb;
  wire [13:0] p3_bit_slice_38197_comb;
  wire [15:0] p3_smul_38199_comb;
  wire [15:0] p3_sub_38200_comb;
  wire [13:0] p3_bit_slice_38201_comb;
  wire [15:0] p3_smul_38203_comb;
  wire [15:0] p3_sub_38204_comb;
  wire [13:0] p3_bit_slice_38205_comb;
  wire [15:0] p3_smul_38207_comb;
  wire [15:0] p3_sub_38208_comb;
  wire [13:0] p3_bit_slice_38209_comb;
  wire [15:0] p3_smul_38211_comb;
  wire [15:0] p3_sub_38212_comb;
  wire [13:0] p3_bit_slice_38213_comb;
  wire [15:0] p3_smul_38215_comb;
  wire [48:0] p3_smul_38217_comb;
  wire [15:0] p3_smul_38218_comb;
  wire [48:0] p3_smul_38220_comb;
  wire [15:0] p3_smul_38221_comb;
  wire [48:0] p3_smul_38223_comb;
  wire [15:0] p3_smul_38224_comb;
  wire [48:0] p3_smul_38226_comb;
  wire [15:0] p3_smul_38227_comb;
  wire [48:0] p3_smul_38229_comb;
  wire [15:0] p3_smul_38230_comb;
  wire [48:0] p3_smul_38232_comb;
  wire [15:0] p3_smul_38233_comb;
  wire [48:0] p3_smul_38235_comb;
  wire [15:0] p3_smul_38236_comb;
  wire [48:0] p3_smul_38238_comb;
  wire [15:0] p3_smul_38239_comb;
  wire [48:0] p3_smul_38241_comb;
  wire [15:0] p3_smul_38242_comb;
  wire [48:0] p3_smul_38244_comb;
  wire [15:0] p3_smul_38245_comb;
  wire [48:0] p3_smul_38247_comb;
  wire [15:0] p3_smul_38248_comb;
  wire [48:0] p3_smul_38250_comb;
  wire [15:0] p3_smul_38251_comb;
  wire [48:0] p3_smul_38253_comb;
  wire [15:0] p3_smul_38254_comb;
  wire [48:0] p3_smul_38256_comb;
  wire [15:0] p3_smul_38257_comb;
  wire [48:0] p3_smul_38259_comb;
  wire [15:0] p3_smul_38260_comb;
  wire [48:0] p3_smul_38262_comb;
  wire [15:0] p3_smul_38263_comb;
  wire [15:0] p3_sub_38264_comb;
  wire [13:0] p3_bit_slice_38265_comb;
  wire [15:0] p3_smul_38267_comb;
  wire [15:0] p3_sub_38268_comb;
  wire [13:0] p3_bit_slice_38269_comb;
  wire [15:0] p3_smul_38271_comb;
  wire [15:0] p3_sub_38272_comb;
  wire [13:0] p3_bit_slice_38273_comb;
  wire [15:0] p3_smul_38275_comb;
  wire [15:0] p3_sub_38276_comb;
  wire [13:0] p3_bit_slice_38277_comb;
  wire [15:0] p3_smul_38279_comb;
  wire [15:0] p3_sub_38280_comb;
  wire [13:0] p3_bit_slice_38281_comb;
  wire [15:0] p3_smul_38283_comb;
  wire [15:0] p3_sub_38284_comb;
  wire [13:0] p3_bit_slice_38285_comb;
  wire [15:0] p3_smul_38287_comb;
  wire [15:0] p3_sub_38288_comb;
  wire [13:0] p3_bit_slice_38289_comb;
  wire [15:0] p3_smul_38291_comb;
  wire [15:0] p3_sub_38292_comb;
  wire [13:0] p3_bit_slice_38293_comb;
  wire [47:0] p3_smul_38329_comb;
  wire [47:0] p3_smul_38332_comb;
  wire [47:0] p3_smul_38335_comb;
  wire [47:0] p3_smul_38338_comb;
  wire [47:0] p3_smul_38341_comb;
  wire [47:0] p3_smul_38344_comb;
  wire [47:0] p3_smul_38347_comb;
  wire [47:0] p3_smul_38350_comb;
  wire [47:0] p3_smul_38353_comb;
  wire [47:0] p3_smul_38356_comb;
  wire [47:0] p3_smul_38359_comb;
  wire [47:0] p3_smul_38362_comb;
  wire [47:0] p3_smul_38365_comb;
  wire [47:0] p3_smul_38368_comb;
  wire [47:0] p3_smul_38371_comb;
  wire [47:0] p3_smul_38374_comb;
  wire [47:0] p3_smul_38441_comb;
  wire [47:0] p3_smul_38444_comb;
  wire [47:0] p3_smul_38447_comb;
  wire [47:0] p3_smul_38450_comb;
  wire [47:0] p3_smul_38453_comb;
  wire [47:0] p3_smul_38456_comb;
  wire [47:0] p3_smul_38459_comb;
  wire [47:0] p3_smul_38462_comb;
  wire [47:0] p3_smul_38464_comb;
  wire [47:0] p3_smul_38466_comb;
  wire [47:0] p3_smul_38468_comb;
  wire [47:0] p3_smul_38470_comb;
  wire [47:0] p3_smul_38472_comb;
  wire [47:0] p3_smul_38474_comb;
  wire [47:0] p3_smul_38476_comb;
  wire [47:0] p3_smul_38478_comb;
  wire [15:0] p3_add_38543_comb;
  wire [15:0] p3_add_38544_comb;
  wire [15:0] p3_add_38545_comb;
  wire [15:0] p3_add_38546_comb;
  wire [15:0] p3_add_38547_comb;
  wire [15:0] p3_add_38548_comb;
  wire [15:0] p3_add_38549_comb;
  wire [15:0] p3_add_38550_comb;
  wire [15:0] p3_add_38551_comb;
  wire [15:0] p3_add_38552_comb;
  wire [15:0] p3_add_38553_comb;
  wire [15:0] p3_add_38554_comb;
  wire [15:0] p3_add_38555_comb;
  wire [15:0] p3_add_38556_comb;
  wire [15:0] p3_add_38557_comb;
  wire [15:0] p3_add_38558_comb;
  wire [15:0] p3_smul_38295_comb;
  wire [15:0] p3_sub_38296_comb;
  wire [13:0] p3_bit_slice_38297_comb;
  wire [15:0] p3_smul_38299_comb;
  wire [15:0] p3_sub_38300_comb;
  wire [13:0] p3_bit_slice_38301_comb;
  wire [15:0] p3_smul_38303_comb;
  wire [15:0] p3_sub_38304_comb;
  wire [13:0] p3_bit_slice_38305_comb;
  wire [15:0] p3_smul_38307_comb;
  wire [15:0] p3_sub_38308_comb;
  wire [13:0] p3_bit_slice_38309_comb;
  wire [15:0] p3_smul_38311_comb;
  wire [15:0] p3_sub_38312_comb;
  wire [13:0] p3_bit_slice_38313_comb;
  wire [15:0] p3_smul_38315_comb;
  wire [15:0] p3_sub_38316_comb;
  wire [13:0] p3_bit_slice_38317_comb;
  wire [15:0] p3_smul_38319_comb;
  wire [15:0] p3_sub_38320_comb;
  wire [13:0] p3_bit_slice_38321_comb;
  wire [15:0] p3_smul_38323_comb;
  wire [15:0] p3_sub_38324_comb;
  wire [13:0] p3_bit_slice_38325_comb;
  wire [15:0] p3_smul_38327_comb;
  wire [15:0] p3_smul_38330_comb;
  wire [15:0] p3_smul_38333_comb;
  wire [15:0] p3_smul_38336_comb;
  wire [15:0] p3_smul_38339_comb;
  wire [15:0] p3_smul_38342_comb;
  wire [15:0] p3_smul_38345_comb;
  wire [15:0] p3_smul_38348_comb;
  wire [12:0] p3_bit_slice_38377_comb;
  wire [12:0] p3_bit_slice_38381_comb;
  wire [12:0] p3_bit_slice_38385_comb;
  wire [12:0] p3_bit_slice_38389_comb;
  wire [12:0] p3_bit_slice_38393_comb;
  wire [12:0] p3_bit_slice_38397_comb;
  wire [12:0] p3_bit_slice_38401_comb;
  wire [12:0] p3_bit_slice_38405_comb;
  wire [12:0] p3_bit_slice_38409_comb;
  wire [12:0] p3_bit_slice_38413_comb;
  wire [12:0] p3_bit_slice_38417_comb;
  wire [12:0] p3_bit_slice_38421_comb;
  wire [12:0] p3_bit_slice_38425_comb;
  wire [12:0] p3_bit_slice_38429_comb;
  wire [12:0] p3_bit_slice_38433_comb;
  wire [12:0] p3_bit_slice_38437_comb;
  wire [12:0] p3_bit_slice_38480_comb;
  wire [12:0] p3_bit_slice_38482_comb;
  wire [12:0] p3_bit_slice_38484_comb;
  wire [12:0] p3_bit_slice_38486_comb;
  wire [12:0] p3_bit_slice_38488_comb;
  wire [12:0] p3_bit_slice_38490_comb;
  wire [12:0] p3_bit_slice_38492_comb;
  wire [12:0] p3_bit_slice_38494_comb;
  wire [12:0] p3_bit_slice_38496_comb;
  wire [12:0] p3_bit_slice_38498_comb;
  wire [12:0] p3_bit_slice_38500_comb;
  wire [12:0] p3_bit_slice_38502_comb;
  wire [12:0] p3_bit_slice_38504_comb;
  wire [12:0] p3_bit_slice_38506_comb;
  wire [12:0] p3_bit_slice_38508_comb;
  wire [12:0] p3_bit_slice_38510_comb;
  wire [15:0] p3_add_38559_comb;
  wire [15:0] p3_add_38560_comb;
  wire [15:0] p3_add_38561_comb;
  wire [15:0] p3_add_38562_comb;
  wire [15:0] p3_add_38563_comb;
  wire [15:0] p3_add_38564_comb;
  wire [15:0] p3_add_38565_comb;
  wire [15:0] p3_add_38566_comb;
  wire [15:0] p3_add_38567_comb;
  wire [15:0] p3_add_38568_comb;
  wire [15:0] p3_add_38569_comb;
  wire [15:0] p3_add_38570_comb;
  wire [15:0] p3_add_38571_comb;
  wire [15:0] p3_add_38572_comb;
  wire [15:0] p3_add_38573_comb;
  wire [15:0] p3_add_38574_comb;
  wire [15:0] p3_add_38575_comb;
  wire [15:0] p3_add_38576_comb;
  wire [15:0] p3_add_38577_comb;
  wire [15:0] p3_add_38579_comb;
  wire [15:0] p3_add_38580_comb;
  wire [15:0] p3_add_38581_comb;
  wire [15:0] p3_add_38583_comb;
  wire [15:0] p3_add_38584_comb;
  wire [15:0] p3_add_38585_comb;
  wire [15:0] p3_add_38587_comb;
  wire [15:0] p3_add_38588_comb;
  wire [15:0] p3_add_38589_comb;
  wire [15:0] p3_add_38591_comb;
  wire [15:0] p3_add_38592_comb;
  wire [15:0] p3_add_38593_comb;
  wire [15:0] p3_add_38595_comb;
  wire [15:0] p3_add_38596_comb;
  wire [15:0] p3_add_38597_comb;
  wire [15:0] p3_add_38599_comb;
  wire [15:0] p3_add_38600_comb;
  wire [15:0] p3_add_38601_comb;
  wire [15:0] p3_add_38603_comb;
  wire [15:0] p3_add_38604_comb;
  wire [15:0] p3_add_38605_comb;
  wire [15:0] p3_smul_38351_comb;
  wire [15:0] p3_smul_38354_comb;
  wire [15:0] p3_smul_38357_comb;
  wire [15:0] p3_smul_38360_comb;
  wire [15:0] p3_smul_38363_comb;
  wire [15:0] p3_smul_38366_comb;
  wire [15:0] p3_smul_38369_comb;
  wire [15:0] p3_smul_38372_comb;
  wire [15:0] p3_smul_38375_comb;
  wire [15:0] p3_sub_38376_comb;
  wire [15:0] p3_smul_38379_comb;
  wire [15:0] p3_sub_38380_comb;
  wire [15:0] p3_smul_38383_comb;
  wire [15:0] p3_sub_38384_comb;
  wire [15:0] p3_smul_38387_comb;
  wire [15:0] p3_sub_38388_comb;
  wire [15:0] p3_smul_38391_comb;
  wire [15:0] p3_sub_38392_comb;
  wire [15:0] p3_smul_38395_comb;
  wire [15:0] p3_sub_38396_comb;
  wire [15:0] p3_smul_38399_comb;
  wire [15:0] p3_sub_38400_comb;
  wire [15:0] p3_smul_38403_comb;
  wire [15:0] p3_sub_38404_comb;
  wire [15:0] p3_add_38607_comb;
  wire [15:0] p3_add_38608_comb;
  wire [15:0] p3_add_38609_comb;
  wire [15:0] p3_add_38610_comb;
  wire [15:0] p3_add_38611_comb;
  wire [15:0] p3_add_38612_comb;
  wire [15:0] p3_add_38613_comb;
  wire [15:0] p3_add_38614_comb;
  wire [15:0] p3_add_38615_comb;
  wire [15:0] p3_add_38616_comb;
  wire [15:0] p3_add_38617_comb;
  wire [15:0] p3_add_38618_comb;
  wire [15:0] p3_add_38619_comb;
  wire [15:0] p3_add_38620_comb;
  wire [15:0] p3_add_38621_comb;
  wire [15:0] p3_add_38622_comb;
  wire [15:0] p3_add_38623_comb;
  wire [15:0] p3_add_38624_comb;
  wire [15:0] p3_add_38625_comb;
  wire [15:0] p3_add_38626_comb;
  wire [15:0] p3_add_38627_comb;
  wire [15:0] p3_add_38628_comb;
  wire [15:0] p3_add_38629_comb;
  wire [15:0] p3_add_38630_comb;
  wire [15:0] p3_add_38631_comb;
  wire [15:0] p3_add_38632_comb;
  wire [15:0] p3_add_38633_comb;
  wire [15:0] p3_add_38634_comb;
  wire [15:0] p3_add_38635_comb;
  wire [15:0] p3_add_38636_comb;
  wire [15:0] p3_add_38637_comb;
  wire [15:0] p3_add_38638_comb;
  wire [15:0] p3_add_38639_comb;
  wire [15:0] p3_add_38640_comb;
  wire [15:0] p3_add_38641_comb;
  wire [15:0] p3_add_38642_comb;
  wire [15:0] p3_add_38643_comb;
  wire [15:0] p3_add_38644_comb;
  wire [15:0] p3_add_38645_comb;
  wire [15:0] p3_add_38646_comb;
  wire [15:0] p3_add_38647_comb;
  wire [15:0] p3_add_38648_comb;
  wire [15:0] p3_add_38649_comb;
  wire [15:0] p3_add_38650_comb;
  wire [15:0] p3_add_38651_comb;
  wire [15:0] p3_add_38652_comb;
  wire [15:0] p3_add_38653_comb;
  wire [15:0] p3_add_38654_comb;
  wire [15:0] p3_smul_38407_comb;
  wire [15:0] p3_sub_38408_comb;
  wire [15:0] p3_smul_38411_comb;
  wire [15:0] p3_sub_38412_comb;
  wire [15:0] p3_smul_38415_comb;
  wire [15:0] p3_sub_38416_comb;
  wire [15:0] p3_smul_38419_comb;
  wire [15:0] p3_sub_38420_comb;
  wire [15:0] p3_smul_38423_comb;
  wire [15:0] p3_sub_38424_comb;
  wire [15:0] p3_smul_38427_comb;
  wire [15:0] p3_sub_38428_comb;
  wire [15:0] p3_smul_38431_comb;
  wire [15:0] p3_sub_38432_comb;
  wire [15:0] p3_smul_38435_comb;
  wire [15:0] p3_sub_38436_comb;
  wire [15:0] p3_smul_38439_comb;
  wire [15:0] p3_smul_38442_comb;
  wire [15:0] p3_smul_38445_comb;
  wire [15:0] p3_smul_38448_comb;
  wire [15:0] p3_smul_38451_comb;
  wire [15:0] p3_smul_38454_comb;
  wire [15:0] p3_smul_38457_comb;
  wire [15:0] p3_smul_38460_comb;
  wire [15:0] p3_sub_38479_comb;
  wire [15:0] p3_sub_38481_comb;
  wire [15:0] p3_sub_38483_comb;
  wire [15:0] p3_sub_38485_comb;
  wire [15:0] p3_sub_38487_comb;
  wire [15:0] p3_sub_38489_comb;
  wire [15:0] p3_sub_38491_comb;
  wire [15:0] p3_sub_38493_comb;
  wire [15:0] p3_sub_38495_comb;
  wire [15:0] p3_sub_38497_comb;
  wire [15:0] p3_sub_38499_comb;
  wire [15:0] p3_sub_38501_comb;
  wire [15:0] p3_sub_38503_comb;
  wire [15:0] p3_sub_38505_comb;
  wire [15:0] p3_sub_38507_comb;
  wire [15:0] p3_sub_38509_comb;
  wire [15:0] p3_sub_38527_comb;
  wire [15:0] p3_sub_38528_comb;
  wire [15:0] p3_sub_38529_comb;
  wire [15:0] p3_sub_38530_comb;
  wire [15:0] p3_sub_38531_comb;
  wire [15:0] p3_sub_38532_comb;
  wire [15:0] p3_sub_38533_comb;
  wire [15:0] p3_sub_38534_comb;
  wire [15:0] p3_sub_38535_comb;
  wire [15:0] p3_sub_38536_comb;
  wire [15:0] p3_sub_38537_comb;
  wire [15:0] p3_sub_38538_comb;
  wire [15:0] p3_sub_38539_comb;
  wire [15:0] p3_sub_38540_comb;
  wire [15:0] p3_sub_38541_comb;
  wire [15:0] p3_sub_38542_comb;
  wire [15:0] p3_add_38578_comb;
  wire [15:0] p3_add_38582_comb;
  wire [15:0] p3_add_38586_comb;
  wire [15:0] p3_add_38590_comb;
  wire [15:0] p3_add_38594_comb;
  wire [15:0] p3_add_38598_comb;
  wire [15:0] p3_add_38602_comb;
  wire [15:0] p3_add_38606_comb;
  wire [15:0] p3_add_38655_comb;
  wire [15:0] p3_add_38656_comb;
  wire [15:0] p3_add_38657_comb;
  wire [15:0] p3_add_38658_comb;
  wire [15:0] p3_add_38659_comb;
  wire [15:0] p3_add_38660_comb;
  wire [15:0] p3_add_38661_comb;
  wire [15:0] p3_add_38662_comb;
  wire [15:0] p3_add_38663_comb;
  wire [15:0] p3_add_38664_comb;
  wire [15:0] p3_add_38665_comb;
  wire [15:0] p3_add_38666_comb;
  wire [15:0] p3_add_38667_comb;
  wire [15:0] p3_add_38668_comb;
  wire [15:0] p3_add_38669_comb;
  wire [15:0] p3_add_38670_comb;
  wire [15:0] p3_add_38671_comb;
  wire [15:0] p3_add_38672_comb;
  wire [15:0] p3_add_38673_comb;
  wire [15:0] p3_add_38674_comb;
  wire [15:0] p3_add_38675_comb;
  wire [15:0] p3_add_38676_comb;
  wire [15:0] p3_add_38677_comb;
  wire [15:0] p3_add_38678_comb;
  assign p3_smul_38023_comb = smul16b_16b_x_16b(p2_smul_37159, p2_sub_37160);
  assign p3_smul_38025_comb = smul16b_16b_x_16b(p2_smul_37164, p2_sub_37165);
  assign p3_smul_38027_comb = smul16b_16b_x_16b(p2_smul_37169, p2_sub_37170);
  assign p3_smul_38029_comb = smul16b_16b_x_16b(p2_smul_37174, p2_sub_37175);
  assign p3_smul_38031_comb = smul16b_16b_x_16b(p2_smul_37179, p2_sub_37180);
  assign p3_smul_38033_comb = smul16b_16b_x_16b(p2_smul_37184, p2_sub_37185);
  assign p3_smul_38035_comb = smul16b_16b_x_16b(p2_smul_37189, p2_sub_37190);
  assign p3_smul_38037_comb = smul16b_16b_x_16b(p2_smul_37194, p2_sub_37195);
  assign p3_smul_38039_comb = smul16b_16b_x_16b(p2_smul_37199, p2_sub_37200);
  assign p3_smul_38040_comb = smul16b_16b_x_16b(p2_smul_37204, p2_sub_37205);
  assign p3_smul_38041_comb = smul16b_16b_x_16b(p2_smul_37209, p2_sub_37210);
  assign p3_smul_38042_comb = smul16b_16b_x_16b(p2_smul_37214, p2_sub_37215);
  assign p3_smul_38043_comb = smul16b_16b_x_16b(p2_smul_37219, p2_sub_37220);
  assign p3_smul_38044_comb = smul16b_16b_x_16b(p2_smul_37224, p2_sub_37225);
  assign p3_smul_38045_comb = smul16b_16b_x_16b(p2_smul_37229, p2_sub_37230);
  assign p3_smul_38046_comb = smul16b_16b_x_16b(p2_smul_37234, p2_sub_37235);
  assign p3_smul_38047_comb = smul16b_16b_x_16b(p3_smul_38023_comb, p2_sub_37239);
  assign p3_smul_38048_comb = smul47b_16b_x_31b(p2_neg_36551, 31'h2e8b_a2e9);
  assign p3_smul_38049_comb = smul16b_16b_x_16b(p3_smul_38025_comb, p2_sub_37242);
  assign p3_smul_38050_comb = smul47b_16b_x_31b(p2_neg_36552, 31'h2e8b_a2e9);
  assign p3_smul_38051_comb = smul16b_16b_x_16b(p3_smul_38027_comb, p2_sub_37245);
  assign p3_smul_38052_comb = smul47b_16b_x_31b(p2_neg_36553, 31'h2e8b_a2e9);
  assign p3_smul_38053_comb = smul16b_16b_x_16b(p3_smul_38029_comb, p2_sub_37248);
  assign p3_smul_38054_comb = smul47b_16b_x_31b(p2_neg_36554, 31'h2e8b_a2e9);
  assign p3_smul_38055_comb = smul16b_16b_x_16b(p3_smul_38031_comb, p2_sub_37251);
  assign p3_smul_38056_comb = smul47b_16b_x_31b(p2_neg_36555, 31'h2e8b_a2e9);
  assign p3_smul_38057_comb = smul16b_16b_x_16b(p3_smul_38033_comb, p2_sub_37254);
  assign p3_smul_38058_comb = smul47b_16b_x_31b(p2_neg_36556, 31'h2e8b_a2e9);
  assign p3_smul_38059_comb = smul16b_16b_x_16b(p3_smul_38035_comb, p2_sub_37257);
  assign p3_smul_38060_comb = smul47b_16b_x_31b(p2_neg_36557, 31'h2e8b_a2e9);
  assign p3_smul_38061_comb = smul16b_16b_x_16b(p3_smul_38037_comb, p2_sub_37260);
  assign p3_smul_38062_comb = smul47b_16b_x_31b(p2_neg_36558, 31'h2e8b_a2e9);
  assign p3_smul_38063_comb = smul16b_16b_x_16b(p3_smul_38039_comb, p2_bit_slice_37263);
  assign p3_smul_38065_comb = smul16b_16b_x_16b(p3_smul_38040_comb, p2_bit_slice_37266);
  assign p3_smul_38067_comb = smul16b_16b_x_16b(p3_smul_38041_comb, p2_bit_slice_37269);
  assign p3_smul_38069_comb = smul16b_16b_x_16b(p3_smul_38042_comb, p2_bit_slice_37272);
  assign p3_smul_38071_comb = smul16b_16b_x_16b(p3_smul_38043_comb, p2_bit_slice_37275);
  assign p3_smul_38073_comb = smul16b_16b_x_16b(p3_smul_38044_comb, p2_bit_slice_37278);
  assign p3_smul_38075_comb = smul16b_16b_x_16b(p3_smul_38045_comb, p2_bit_slice_37281);
  assign p3_smul_38077_comb = smul16b_16b_x_16b(p3_smul_38046_comb, p2_bit_slice_37284);
  assign p3_smul_38079_comb = smul16b_16b_x_16b(p3_smul_38047_comb, p2_bit_slice_37287);
  assign p3_bit_slice_38080_comb = p3_smul_38048_comb[46:33];
  assign p3_smul_38082_comb = smul16b_16b_x_16b(p3_smul_38049_comb, p2_bit_slice_37289);
  assign p3_bit_slice_38083_comb = p3_smul_38050_comb[46:33];
  assign p3_smul_38085_comb = smul16b_16b_x_16b(p3_smul_38051_comb, p2_bit_slice_37291);
  assign p3_bit_slice_38086_comb = p3_smul_38052_comb[46:33];
  assign p3_smul_38088_comb = smul16b_16b_x_16b(p3_smul_38053_comb, p2_bit_slice_37293);
  assign p3_bit_slice_38089_comb = p3_smul_38054_comb[46:33];
  assign p3_smul_38091_comb = smul16b_16b_x_16b(p3_smul_38055_comb, p2_bit_slice_37295);
  assign p3_bit_slice_38092_comb = p3_smul_38056_comb[46:33];
  assign p3_smul_38094_comb = smul16b_16b_x_16b(p3_smul_38057_comb, p2_bit_slice_37297);
  assign p3_bit_slice_38095_comb = p3_smul_38058_comb[46:33];
  assign p3_smul_38097_comb = smul16b_16b_x_16b(p3_smul_38059_comb, p2_bit_slice_37299);
  assign p3_bit_slice_38098_comb = p3_smul_38060_comb[46:33];
  assign p3_smul_38100_comb = smul16b_16b_x_16b(p3_smul_38061_comb, p2_bit_slice_37301);
  assign p3_bit_slice_38101_comb = p3_smul_38062_comb[46:33];
  assign p3_smul_38103_comb = smul16b_16b_x_16b(p3_smul_38063_comb, p2_sub_37303);
  assign p3_smul_38105_comb = smul48b_16b_x_32b(p2_neg_36543, 32'h4ec4_ec4f);
  assign p3_smul_38106_comb = smul16b_16b_x_16b(p3_smul_38065_comb, p2_sub_37306);
  assign p3_smul_38108_comb = smul48b_16b_x_32b(p2_neg_36544, 32'h4ec4_ec4f);
  assign p3_smul_38109_comb = smul16b_16b_x_16b(p3_smul_38067_comb, p2_sub_37309);
  assign p3_smul_38111_comb = smul48b_16b_x_32b(p2_neg_36545, 32'h4ec4_ec4f);
  assign p3_smul_38112_comb = smul16b_16b_x_16b(p3_smul_38069_comb, p2_sub_37312);
  assign p3_smul_38114_comb = smul48b_16b_x_32b(p2_neg_36546, 32'h4ec4_ec4f);
  assign p3_smul_38115_comb = smul16b_16b_x_16b(p3_smul_38071_comb, p2_sub_37315);
  assign p3_smul_38117_comb = smul48b_16b_x_32b(p2_neg_36547, 32'h4ec4_ec4f);
  assign p3_smul_38118_comb = smul16b_16b_x_16b(p3_smul_38073_comb, p2_sub_37318);
  assign p3_smul_38120_comb = smul48b_16b_x_32b(p2_neg_36548, 32'h4ec4_ec4f);
  assign p3_smul_38121_comb = smul16b_16b_x_16b(p3_smul_38075_comb, p2_sub_37321);
  assign p3_smul_38123_comb = smul48b_16b_x_32b(p2_neg_36549, 32'h4ec4_ec4f);
  assign p3_smul_38124_comb = smul16b_16b_x_16b(p3_smul_38077_comb, p2_sub_37324);
  assign p3_smul_38126_comb = smul48b_16b_x_32b(p2_neg_36550, 32'h4ec4_ec4f);
  assign p3_smul_38127_comb = smul16b_16b_x_16b(p3_smul_38079_comb, p2_sub_37327);
  assign p3_smul_38129_comb = smul48b_16b_x_32b(p2_neg_36551, 32'h4ec4_ec4f);
  assign p3_smul_38130_comb = smul16b_16b_x_16b(p3_smul_38082_comb, p2_sub_37329);
  assign p3_smul_38132_comb = smul48b_16b_x_32b(p2_neg_36552, 32'h4ec4_ec4f);
  assign p3_smul_38133_comb = smul16b_16b_x_16b(p3_smul_38085_comb, p2_sub_37331);
  assign p3_smul_38135_comb = smul48b_16b_x_32b(p2_neg_36553, 32'h4ec4_ec4f);
  assign p3_smul_38136_comb = smul16b_16b_x_16b(p3_smul_38088_comb, p2_sub_37333);
  assign p3_smul_38138_comb = smul48b_16b_x_32b(p2_neg_36554, 32'h4ec4_ec4f);
  assign p3_smul_38139_comb = smul16b_16b_x_16b(p3_smul_38091_comb, p2_sub_37335);
  assign p3_smul_38141_comb = smul48b_16b_x_32b(p2_neg_36555, 32'h4ec4_ec4f);
  assign p3_smul_38142_comb = smul16b_16b_x_16b(p3_smul_38094_comb, p2_sub_37337);
  assign p3_smul_38144_comb = smul48b_16b_x_32b(p2_neg_36556, 32'h4ec4_ec4f);
  assign p3_smul_38145_comb = smul16b_16b_x_16b(p3_smul_38097_comb, p2_sub_37339);
  assign p3_smul_38147_comb = smul48b_16b_x_32b(p2_neg_36557, 32'h4ec4_ec4f);
  assign p3_smul_38148_comb = smul16b_16b_x_16b(p3_smul_38100_comb, p2_sub_37341);
  assign p3_smul_38150_comb = smul48b_16b_x_32b(p2_neg_36558, 32'h4ec4_ec4f);
  assign p3_smul_38151_comb = smul16b_16b_x_16b(p3_smul_38103_comb, p2_sub_37343);
  assign p3_sub_38152_comb = {{2{p2_bit_slice_37305[13]}}, p2_bit_slice_37305} - p2_sign_ext_36769;
  assign p3_bit_slice_38153_comb = p3_smul_38105_comb[47:34];
  assign p3_smul_38155_comb = smul16b_16b_x_16b(p3_smul_38106_comb, p2_sub_37344);
  assign p3_sub_38156_comb = {{2{p2_bit_slice_37308[13]}}, p2_bit_slice_37308} - p2_sign_ext_36774;
  assign p3_bit_slice_38157_comb = p3_smul_38108_comb[47:34];
  assign p3_smul_38159_comb = smul16b_16b_x_16b(p3_smul_38109_comb, p2_sub_37345);
  assign p3_sub_38160_comb = {{2{p2_bit_slice_37311[13]}}, p2_bit_slice_37311} - p2_sign_ext_36779;
  assign p3_bit_slice_38161_comb = p3_smul_38111_comb[47:34];
  assign p3_smul_38163_comb = smul16b_16b_x_16b(p3_smul_38112_comb, p2_sub_37346);
  assign p3_sub_38164_comb = {{2{p2_bit_slice_37314[13]}}, p2_bit_slice_37314} - p2_sign_ext_36784;
  assign p3_bit_slice_38165_comb = p3_smul_38114_comb[47:34];
  assign p3_smul_38167_comb = smul16b_16b_x_16b(p3_smul_38115_comb, p2_sub_37347);
  assign p3_sub_38168_comb = {{2{p2_bit_slice_37317[13]}}, p2_bit_slice_37317} - p2_sign_ext_36789;
  assign p3_bit_slice_38169_comb = p3_smul_38117_comb[47:34];
  assign p3_smul_38171_comb = smul16b_16b_x_16b(p3_smul_38118_comb, p2_sub_37348);
  assign p3_sub_38172_comb = {{2{p2_bit_slice_37320[13]}}, p2_bit_slice_37320} - p2_sign_ext_36794;
  assign p3_bit_slice_38173_comb = p3_smul_38120_comb[47:34];
  assign p3_smul_38175_comb = smul16b_16b_x_16b(p3_smul_38121_comb, p2_sub_37349);
  assign p3_sub_38176_comb = {{2{p2_bit_slice_37323[13]}}, p2_bit_slice_37323} - p2_sign_ext_36799;
  assign p3_bit_slice_38177_comb = p3_smul_38123_comb[47:34];
  assign p3_smul_38179_comb = smul16b_16b_x_16b(p3_smul_38124_comb, p2_sub_37350);
  assign p3_sub_38180_comb = {{2{p2_bit_slice_37326[13]}}, p2_bit_slice_37326} - p2_sign_ext_36804;
  assign p3_bit_slice_38181_comb = p3_smul_38126_comb[47:34];
  assign p3_smul_38183_comb = smul16b_16b_x_16b(p3_smul_38127_comb, p2_sub_37351);
  assign p3_sub_38184_comb = {{2{p3_bit_slice_38080_comb[13]}}, p3_bit_slice_38080_comb} - p2_sign_ext_36809;
  assign p3_bit_slice_38185_comb = p3_smul_38129_comb[47:34];
  assign p3_smul_38187_comb = smul16b_16b_x_16b(p3_smul_38130_comb, p2_sub_37352);
  assign p3_sub_38188_comb = {{2{p3_bit_slice_38083_comb[13]}}, p3_bit_slice_38083_comb} - p2_sign_ext_36814;
  assign p3_bit_slice_38189_comb = p3_smul_38132_comb[47:34];
  assign p3_smul_38191_comb = smul16b_16b_x_16b(p3_smul_38133_comb, p2_sub_37353);
  assign p3_sub_38192_comb = {{2{p3_bit_slice_38086_comb[13]}}, p3_bit_slice_38086_comb} - p2_sign_ext_36819;
  assign p3_bit_slice_38193_comb = p3_smul_38135_comb[47:34];
  assign p3_smul_38195_comb = smul16b_16b_x_16b(p3_smul_38136_comb, p2_sub_37354);
  assign p3_sub_38196_comb = {{2{p3_bit_slice_38089_comb[13]}}, p3_bit_slice_38089_comb} - p2_sign_ext_36824;
  assign p3_bit_slice_38197_comb = p3_smul_38138_comb[47:34];
  assign p3_smul_38199_comb = smul16b_16b_x_16b(p3_smul_38139_comb, p2_sub_37355);
  assign p3_sub_38200_comb = {{2{p3_bit_slice_38092_comb[13]}}, p3_bit_slice_38092_comb} - p2_sign_ext_36829;
  assign p3_bit_slice_38201_comb = p3_smul_38141_comb[47:34];
  assign p3_smul_38203_comb = smul16b_16b_x_16b(p3_smul_38142_comb, p2_sub_37356);
  assign p3_sub_38204_comb = {{2{p3_bit_slice_38095_comb[13]}}, p3_bit_slice_38095_comb} - p2_sign_ext_36834;
  assign p3_bit_slice_38205_comb = p3_smul_38144_comb[47:34];
  assign p3_smul_38207_comb = smul16b_16b_x_16b(p3_smul_38145_comb, p2_sub_37357);
  assign p3_sub_38208_comb = {{2{p3_bit_slice_38098_comb[13]}}, p3_bit_slice_38098_comb} - p2_sign_ext_36839;
  assign p3_bit_slice_38209_comb = p3_smul_38147_comb[47:34];
  assign p3_smul_38211_comb = smul16b_16b_x_16b(p3_smul_38148_comb, p2_sub_37358);
  assign p3_sub_38212_comb = {{2{p3_bit_slice_38101_comb[13]}}, p3_bit_slice_38101_comb} - p2_sign_ext_36844;
  assign p3_bit_slice_38213_comb = p3_smul_38150_comb[47:34];
  assign p3_smul_38215_comb = smul16b_16b_x_16b(p3_smul_38151_comb, p3_sub_38152_comb);
  assign p3_smul_38217_comb = smul49b_16b_x_33b(p2_neg_36543, 33'h0_8888_8889);
  assign p3_smul_38218_comb = smul16b_16b_x_16b(p3_smul_38155_comb, p3_sub_38156_comb);
  assign p3_smul_38220_comb = smul49b_16b_x_33b(p2_neg_36544, 33'h0_8888_8889);
  assign p3_smul_38221_comb = smul16b_16b_x_16b(p3_smul_38159_comb, p3_sub_38160_comb);
  assign p3_smul_38223_comb = smul49b_16b_x_33b(p2_neg_36545, 33'h0_8888_8889);
  assign p3_smul_38224_comb = smul16b_16b_x_16b(p3_smul_38163_comb, p3_sub_38164_comb);
  assign p3_smul_38226_comb = smul49b_16b_x_33b(p2_neg_36546, 33'h0_8888_8889);
  assign p3_smul_38227_comb = smul16b_16b_x_16b(p3_smul_38167_comb, p3_sub_38168_comb);
  assign p3_smul_38229_comb = smul49b_16b_x_33b(p2_neg_36547, 33'h0_8888_8889);
  assign p3_smul_38230_comb = smul16b_16b_x_16b(p3_smul_38171_comb, p3_sub_38172_comb);
  assign p3_smul_38232_comb = smul49b_16b_x_33b(p2_neg_36548, 33'h0_8888_8889);
  assign p3_smul_38233_comb = smul16b_16b_x_16b(p3_smul_38175_comb, p3_sub_38176_comb);
  assign p3_smul_38235_comb = smul49b_16b_x_33b(p2_neg_36549, 33'h0_8888_8889);
  assign p3_smul_38236_comb = smul16b_16b_x_16b(p3_smul_38179_comb, p3_sub_38180_comb);
  assign p3_smul_38238_comb = smul49b_16b_x_33b(p2_neg_36550, 33'h0_8888_8889);
  assign p3_smul_38239_comb = smul16b_16b_x_16b(p3_smul_38183_comb, p3_sub_38184_comb);
  assign p3_smul_38241_comb = smul49b_16b_x_33b(p2_neg_36551, 33'h0_8888_8889);
  assign p3_smul_38242_comb = smul16b_16b_x_16b(p3_smul_38187_comb, p3_sub_38188_comb);
  assign p3_smul_38244_comb = smul49b_16b_x_33b(p2_neg_36552, 33'h0_8888_8889);
  assign p3_smul_38245_comb = smul16b_16b_x_16b(p3_smul_38191_comb, p3_sub_38192_comb);
  assign p3_smul_38247_comb = smul49b_16b_x_33b(p2_neg_36553, 33'h0_8888_8889);
  assign p3_smul_38248_comb = smul16b_16b_x_16b(p3_smul_38195_comb, p3_sub_38196_comb);
  assign p3_smul_38250_comb = smul49b_16b_x_33b(p2_neg_36554, 33'h0_8888_8889);
  assign p3_smul_38251_comb = smul16b_16b_x_16b(p3_smul_38199_comb, p3_sub_38200_comb);
  assign p3_smul_38253_comb = smul49b_16b_x_33b(p2_neg_36555, 33'h0_8888_8889);
  assign p3_smul_38254_comb = smul16b_16b_x_16b(p3_smul_38203_comb, p3_sub_38204_comb);
  assign p3_smul_38256_comb = smul49b_16b_x_33b(p2_neg_36556, 33'h0_8888_8889);
  assign p3_smul_38257_comb = smul16b_16b_x_16b(p3_smul_38207_comb, p3_sub_38208_comb);
  assign p3_smul_38259_comb = smul49b_16b_x_33b(p2_neg_36557, 33'h0_8888_8889);
  assign p3_smul_38260_comb = smul16b_16b_x_16b(p3_smul_38211_comb, p3_sub_38212_comb);
  assign p3_smul_38262_comb = smul49b_16b_x_33b(p2_neg_36558, 33'h0_8888_8889);
  assign p3_smul_38263_comb = smul16b_16b_x_16b(p3_smul_38215_comb, p2_sub_37375);
  assign p3_sub_38264_comb = {{2{p3_bit_slice_38153_comb[13]}}, p3_bit_slice_38153_comb} - p2_sign_ext_36769;
  assign p3_bit_slice_38265_comb = p3_smul_38217_comb[48:35];
  assign p3_smul_38267_comb = smul16b_16b_x_16b(p3_smul_38218_comb, p2_sub_37376);
  assign p3_sub_38268_comb = {{2{p3_bit_slice_38157_comb[13]}}, p3_bit_slice_38157_comb} - p2_sign_ext_36774;
  assign p3_bit_slice_38269_comb = p3_smul_38220_comb[48:35];
  assign p3_smul_38271_comb = smul16b_16b_x_16b(p3_smul_38221_comb, p2_sub_37377);
  assign p3_sub_38272_comb = {{2{p3_bit_slice_38161_comb[13]}}, p3_bit_slice_38161_comb} - p2_sign_ext_36779;
  assign p3_bit_slice_38273_comb = p3_smul_38223_comb[48:35];
  assign p3_smul_38275_comb = smul16b_16b_x_16b(p3_smul_38224_comb, p2_sub_37378);
  assign p3_sub_38276_comb = {{2{p3_bit_slice_38165_comb[13]}}, p3_bit_slice_38165_comb} - p2_sign_ext_36784;
  assign p3_bit_slice_38277_comb = p3_smul_38226_comb[48:35];
  assign p3_smul_38279_comb = smul16b_16b_x_16b(p3_smul_38227_comb, p2_sub_37379);
  assign p3_sub_38280_comb = {{2{p3_bit_slice_38169_comb[13]}}, p3_bit_slice_38169_comb} - p2_sign_ext_36789;
  assign p3_bit_slice_38281_comb = p3_smul_38229_comb[48:35];
  assign p3_smul_38283_comb = smul16b_16b_x_16b(p3_smul_38230_comb, p2_sub_37380);
  assign p3_sub_38284_comb = {{2{p3_bit_slice_38173_comb[13]}}, p3_bit_slice_38173_comb} - p2_sign_ext_36794;
  assign p3_bit_slice_38285_comb = p3_smul_38232_comb[48:35];
  assign p3_smul_38287_comb = smul16b_16b_x_16b(p3_smul_38233_comb, p2_sub_37381);
  assign p3_sub_38288_comb = {{2{p3_bit_slice_38177_comb[13]}}, p3_bit_slice_38177_comb} - p2_sign_ext_36799;
  assign p3_bit_slice_38289_comb = p3_smul_38235_comb[48:35];
  assign p3_smul_38291_comb = smul16b_16b_x_16b(p3_smul_38236_comb, p2_sub_37382);
  assign p3_sub_38292_comb = {{2{p3_bit_slice_38181_comb[13]}}, p3_bit_slice_38181_comb} - p2_sign_ext_36804;
  assign p3_bit_slice_38293_comb = p3_smul_38238_comb[48:35];
  assign p3_smul_38329_comb = smul48b_16b_x_32b(p2_neg_36543, 32'h7878_7879);
  assign p3_smul_38332_comb = smul48b_16b_x_32b(p2_neg_36544, 32'h7878_7879);
  assign p3_smul_38335_comb = smul48b_16b_x_32b(p2_neg_36545, 32'h7878_7879);
  assign p3_smul_38338_comb = smul48b_16b_x_32b(p2_neg_36546, 32'h7878_7879);
  assign p3_smul_38341_comb = smul48b_16b_x_32b(p2_neg_36547, 32'h7878_7879);
  assign p3_smul_38344_comb = smul48b_16b_x_32b(p2_neg_36548, 32'h7878_7879);
  assign p3_smul_38347_comb = smul48b_16b_x_32b(p2_neg_36549, 32'h7878_7879);
  assign p3_smul_38350_comb = smul48b_16b_x_32b(p2_neg_36550, 32'h7878_7879);
  assign p3_smul_38353_comb = smul48b_16b_x_32b(p2_neg_36551, 32'h7878_7879);
  assign p3_smul_38356_comb = smul48b_16b_x_32b(p2_neg_36552, 32'h7878_7879);
  assign p3_smul_38359_comb = smul48b_16b_x_32b(p2_neg_36553, 32'h7878_7879);
  assign p3_smul_38362_comb = smul48b_16b_x_32b(p2_neg_36554, 32'h7878_7879);
  assign p3_smul_38365_comb = smul48b_16b_x_32b(p2_neg_36555, 32'h7878_7879);
  assign p3_smul_38368_comb = smul48b_16b_x_32b(p2_neg_36556, 32'h7878_7879);
  assign p3_smul_38371_comb = smul48b_16b_x_32b(p2_neg_36557, 32'h7878_7879);
  assign p3_smul_38374_comb = smul48b_16b_x_32b(p2_neg_36558, 32'h7878_7879);
  assign p3_smul_38441_comb = smul48b_16b_x_32b(p2_neg_36543, 32'h6bca_1af3);
  assign p3_smul_38444_comb = smul48b_16b_x_32b(p2_neg_36544, 32'h6bca_1af3);
  assign p3_smul_38447_comb = smul48b_16b_x_32b(p2_neg_36545, 32'h6bca_1af3);
  assign p3_smul_38450_comb = smul48b_16b_x_32b(p2_neg_36546, 32'h6bca_1af3);
  assign p3_smul_38453_comb = smul48b_16b_x_32b(p2_neg_36547, 32'h6bca_1af3);
  assign p3_smul_38456_comb = smul48b_16b_x_32b(p2_neg_36548, 32'h6bca_1af3);
  assign p3_smul_38459_comb = smul48b_16b_x_32b(p2_neg_36549, 32'h6bca_1af3);
  assign p3_smul_38462_comb = smul48b_16b_x_32b(p2_neg_36550, 32'h6bca_1af3);
  assign p3_smul_38464_comb = smul48b_16b_x_32b(p2_neg_36551, 32'h6bca_1af3);
  assign p3_smul_38466_comb = smul48b_16b_x_32b(p2_neg_36552, 32'h6bca_1af3);
  assign p3_smul_38468_comb = smul48b_16b_x_32b(p2_neg_36553, 32'h6bca_1af3);
  assign p3_smul_38470_comb = smul48b_16b_x_32b(p2_neg_36554, 32'h6bca_1af3);
  assign p3_smul_38472_comb = smul48b_16b_x_32b(p2_neg_36555, 32'h6bca_1af3);
  assign p3_smul_38474_comb = smul48b_16b_x_32b(p2_neg_36556, 32'h6bca_1af3);
  assign p3_smul_38476_comb = smul48b_16b_x_32b(p2_neg_36557, 32'h6bca_1af3);
  assign p3_smul_38478_comb = smul48b_16b_x_32b(p2_neg_36558, 32'h6bca_1af3);
  assign p3_add_38543_comb = p2_smul_37119 + p2_smul_37199;
  assign p3_add_38544_comb = p3_smul_38039_comb + p3_smul_38063_comb;
  assign p3_add_38545_comb = p2_smul_37124 + p2_smul_37204;
  assign p3_add_38546_comb = p3_smul_38040_comb + p3_smul_38065_comb;
  assign p3_add_38547_comb = p2_smul_37129 + p2_smul_37209;
  assign p3_add_38548_comb = p3_smul_38041_comb + p3_smul_38067_comb;
  assign p3_add_38549_comb = p2_smul_37134 + p2_smul_37214;
  assign p3_add_38550_comb = p3_smul_38042_comb + p3_smul_38069_comb;
  assign p3_add_38551_comb = p2_smul_37139 + p2_smul_37219;
  assign p3_add_38552_comb = p3_smul_38043_comb + p3_smul_38071_comb;
  assign p3_add_38553_comb = p2_smul_37144 + p2_smul_37224;
  assign p3_add_38554_comb = p3_smul_38044_comb + p3_smul_38073_comb;
  assign p3_add_38555_comb = p2_smul_37149 + p2_smul_37229;
  assign p3_add_38556_comb = p3_smul_38045_comb + p3_smul_38075_comb;
  assign p3_add_38557_comb = p2_smul_37154 + p2_smul_37234;
  assign p3_add_38558_comb = p3_smul_38046_comb + p3_smul_38077_comb;
  assign p3_smul_38295_comb = smul16b_16b_x_16b(p3_smul_38239_comb, p2_sub_37383);
  assign p3_sub_38296_comb = {{2{p3_bit_slice_38185_comb[13]}}, p3_bit_slice_38185_comb} - p2_sign_ext_36809;
  assign p3_bit_slice_38297_comb = p3_smul_38241_comb[48:35];
  assign p3_smul_38299_comb = smul16b_16b_x_16b(p3_smul_38242_comb, p2_sub_37384);
  assign p3_sub_38300_comb = {{2{p3_bit_slice_38189_comb[13]}}, p3_bit_slice_38189_comb} - p2_sign_ext_36814;
  assign p3_bit_slice_38301_comb = p3_smul_38244_comb[48:35];
  assign p3_smul_38303_comb = smul16b_16b_x_16b(p3_smul_38245_comb, p2_sub_37385);
  assign p3_sub_38304_comb = {{2{p3_bit_slice_38193_comb[13]}}, p3_bit_slice_38193_comb} - p2_sign_ext_36819;
  assign p3_bit_slice_38305_comb = p3_smul_38247_comb[48:35];
  assign p3_smul_38307_comb = smul16b_16b_x_16b(p3_smul_38248_comb, p2_sub_37386);
  assign p3_sub_38308_comb = {{2{p3_bit_slice_38197_comb[13]}}, p3_bit_slice_38197_comb} - p2_sign_ext_36824;
  assign p3_bit_slice_38309_comb = p3_smul_38250_comb[48:35];
  assign p3_smul_38311_comb = smul16b_16b_x_16b(p3_smul_38251_comb, p2_sub_37387);
  assign p3_sub_38312_comb = {{2{p3_bit_slice_38201_comb[13]}}, p3_bit_slice_38201_comb} - p2_sign_ext_36829;
  assign p3_bit_slice_38313_comb = p3_smul_38253_comb[48:35];
  assign p3_smul_38315_comb = smul16b_16b_x_16b(p3_smul_38254_comb, p2_sub_37388);
  assign p3_sub_38316_comb = {{2{p3_bit_slice_38205_comb[13]}}, p3_bit_slice_38205_comb} - p2_sign_ext_36834;
  assign p3_bit_slice_38317_comb = p3_smul_38256_comb[48:35];
  assign p3_smul_38319_comb = smul16b_16b_x_16b(p3_smul_38257_comb, p2_sub_37389);
  assign p3_sub_38320_comb = {{2{p3_bit_slice_38209_comb[13]}}, p3_bit_slice_38209_comb} - p2_sign_ext_36839;
  assign p3_bit_slice_38321_comb = p3_smul_38259_comb[48:35];
  assign p3_smul_38323_comb = smul16b_16b_x_16b(p3_smul_38260_comb, p2_sub_37390);
  assign p3_sub_38324_comb = {{2{p3_bit_slice_38213_comb[13]}}, p3_bit_slice_38213_comb} - p2_sign_ext_36844;
  assign p3_bit_slice_38325_comb = p3_smul_38262_comb[48:35];
  assign p3_smul_38327_comb = smul16b_16b_x_16b(p3_smul_38263_comb, p3_sub_38264_comb);
  assign p3_smul_38330_comb = smul16b_16b_x_16b(p3_smul_38267_comb, p3_sub_38268_comb);
  assign p3_smul_38333_comb = smul16b_16b_x_16b(p3_smul_38271_comb, p3_sub_38272_comb);
  assign p3_smul_38336_comb = smul16b_16b_x_16b(p3_smul_38275_comb, p3_sub_38276_comb);
  assign p3_smul_38339_comb = smul16b_16b_x_16b(p3_smul_38279_comb, p3_sub_38280_comb);
  assign p3_smul_38342_comb = smul16b_16b_x_16b(p3_smul_38283_comb, p3_sub_38284_comb);
  assign p3_smul_38345_comb = smul16b_16b_x_16b(p3_smul_38287_comb, p3_sub_38288_comb);
  assign p3_smul_38348_comb = smul16b_16b_x_16b(p3_smul_38291_comb, p3_sub_38292_comb);
  assign p3_bit_slice_38377_comb = p3_smul_38329_comb[47:35];
  assign p3_bit_slice_38381_comb = p3_smul_38332_comb[47:35];
  assign p3_bit_slice_38385_comb = p3_smul_38335_comb[47:35];
  assign p3_bit_slice_38389_comb = p3_smul_38338_comb[47:35];
  assign p3_bit_slice_38393_comb = p3_smul_38341_comb[47:35];
  assign p3_bit_slice_38397_comb = p3_smul_38344_comb[47:35];
  assign p3_bit_slice_38401_comb = p3_smul_38347_comb[47:35];
  assign p3_bit_slice_38405_comb = p3_smul_38350_comb[47:35];
  assign p3_bit_slice_38409_comb = p3_smul_38353_comb[47:35];
  assign p3_bit_slice_38413_comb = p3_smul_38356_comb[47:35];
  assign p3_bit_slice_38417_comb = p3_smul_38359_comb[47:35];
  assign p3_bit_slice_38421_comb = p3_smul_38362_comb[47:35];
  assign p3_bit_slice_38425_comb = p3_smul_38365_comb[47:35];
  assign p3_bit_slice_38429_comb = p3_smul_38368_comb[47:35];
  assign p3_bit_slice_38433_comb = p3_smul_38371_comb[47:35];
  assign p3_bit_slice_38437_comb = p3_smul_38374_comb[47:35];
  assign p3_bit_slice_38480_comb = p3_smul_38441_comb[47:35];
  assign p3_bit_slice_38482_comb = p3_smul_38444_comb[47:35];
  assign p3_bit_slice_38484_comb = p3_smul_38447_comb[47:35];
  assign p3_bit_slice_38486_comb = p3_smul_38450_comb[47:35];
  assign p3_bit_slice_38488_comb = p3_smul_38453_comb[47:35];
  assign p3_bit_slice_38490_comb = p3_smul_38456_comb[47:35];
  assign p3_bit_slice_38492_comb = p3_smul_38459_comb[47:35];
  assign p3_bit_slice_38494_comb = p3_smul_38462_comb[47:35];
  assign p3_bit_slice_38496_comb = p3_smul_38464_comb[47:35];
  assign p3_bit_slice_38498_comb = p3_smul_38466_comb[47:35];
  assign p3_bit_slice_38500_comb = p3_smul_38468_comb[47:35];
  assign p3_bit_slice_38502_comb = p3_smul_38470_comb[47:35];
  assign p3_bit_slice_38504_comb = p3_smul_38472_comb[47:35];
  assign p3_bit_slice_38506_comb = p3_smul_38474_comb[47:35];
  assign p3_bit_slice_38508_comb = p3_smul_38476_comb[47:35];
  assign p3_bit_slice_38510_comb = p3_smul_38478_comb[47:35];
  assign p3_add_38559_comb = p2_smul_37159 + p3_smul_38023_comb;
  assign p3_add_38560_comb = p3_smul_38047_comb + p3_smul_38079_comb;
  assign p3_add_38561_comb = p2_smul_37164 + p3_smul_38025_comb;
  assign p3_add_38562_comb = p3_smul_38049_comb + p3_smul_38082_comb;
  assign p3_add_38563_comb = p2_smul_37169 + p3_smul_38027_comb;
  assign p3_add_38564_comb = p3_smul_38051_comb + p3_smul_38085_comb;
  assign p3_add_38565_comb = p2_smul_37174 + p3_smul_38029_comb;
  assign p3_add_38566_comb = p3_smul_38053_comb + p3_smul_38088_comb;
  assign p3_add_38567_comb = p2_smul_37179 + p3_smul_38031_comb;
  assign p3_add_38568_comb = p3_smul_38055_comb + p3_smul_38091_comb;
  assign p3_add_38569_comb = p2_smul_37184 + p3_smul_38033_comb;
  assign p3_add_38570_comb = p3_smul_38057_comb + p3_smul_38094_comb;
  assign p3_add_38571_comb = p2_smul_37189 + p3_smul_38035_comb;
  assign p3_add_38572_comb = p3_smul_38059_comb + p3_smul_38097_comb;
  assign p3_add_38573_comb = p2_smul_37194 + p3_smul_38037_comb;
  assign p3_add_38574_comb = p3_smul_38061_comb + p3_smul_38100_comb;
  assign p3_add_38575_comb = p3_add_38543_comb + p3_add_38544_comb;
  assign p3_add_38576_comb = p3_smul_38103_comb + p3_smul_38151_comb;
  assign p3_add_38577_comb = p3_smul_38215_comb + p3_smul_38263_comb;
  assign p3_add_38579_comb = p3_add_38545_comb + p3_add_38546_comb;
  assign p3_add_38580_comb = p3_smul_38106_comb + p3_smul_38155_comb;
  assign p3_add_38581_comb = p3_smul_38218_comb + p3_smul_38267_comb;
  assign p3_add_38583_comb = p3_add_38547_comb + p3_add_38548_comb;
  assign p3_add_38584_comb = p3_smul_38109_comb + p3_smul_38159_comb;
  assign p3_add_38585_comb = p3_smul_38221_comb + p3_smul_38271_comb;
  assign p3_add_38587_comb = p3_add_38549_comb + p3_add_38550_comb;
  assign p3_add_38588_comb = p3_smul_38112_comb + p3_smul_38163_comb;
  assign p3_add_38589_comb = p3_smul_38224_comb + p3_smul_38275_comb;
  assign p3_add_38591_comb = p3_add_38551_comb + p3_add_38552_comb;
  assign p3_add_38592_comb = p3_smul_38115_comb + p3_smul_38167_comb;
  assign p3_add_38593_comb = p3_smul_38227_comb + p3_smul_38279_comb;
  assign p3_add_38595_comb = p3_add_38553_comb + p3_add_38554_comb;
  assign p3_add_38596_comb = p3_smul_38118_comb + p3_smul_38171_comb;
  assign p3_add_38597_comb = p3_smul_38230_comb + p3_smul_38283_comb;
  assign p3_add_38599_comb = p3_add_38555_comb + p3_add_38556_comb;
  assign p3_add_38600_comb = p3_smul_38121_comb + p3_smul_38175_comb;
  assign p3_add_38601_comb = p3_smul_38233_comb + p3_smul_38287_comb;
  assign p3_add_38603_comb = p3_add_38557_comb + p3_add_38558_comb;
  assign p3_add_38604_comb = p3_smul_38124_comb + p3_smul_38179_comb;
  assign p3_add_38605_comb = p3_smul_38236_comb + p3_smul_38291_comb;
  assign p3_smul_38351_comb = smul16b_16b_x_16b(p3_smul_38295_comb, p3_sub_38296_comb);
  assign p3_smul_38354_comb = smul16b_16b_x_16b(p3_smul_38299_comb, p3_sub_38300_comb);
  assign p3_smul_38357_comb = smul16b_16b_x_16b(p3_smul_38303_comb, p3_sub_38304_comb);
  assign p3_smul_38360_comb = smul16b_16b_x_16b(p3_smul_38307_comb, p3_sub_38308_comb);
  assign p3_smul_38363_comb = smul16b_16b_x_16b(p3_smul_38311_comb, p3_sub_38312_comb);
  assign p3_smul_38366_comb = smul16b_16b_x_16b(p3_smul_38315_comb, p3_sub_38316_comb);
  assign p3_smul_38369_comb = smul16b_16b_x_16b(p3_smul_38319_comb, p3_sub_38320_comb);
  assign p3_smul_38372_comb = smul16b_16b_x_16b(p3_smul_38323_comb, p3_sub_38324_comb);
  assign p3_smul_38375_comb = smul16b_16b_x_16b(p3_smul_38327_comb, p2_sub_37439);
  assign p3_sub_38376_comb = {{2{p3_bit_slice_38265_comb[13]}}, p3_bit_slice_38265_comb} - p2_sign_ext_36769;
  assign p3_smul_38379_comb = smul16b_16b_x_16b(p3_smul_38330_comb, p2_sub_37441);
  assign p3_sub_38380_comb = {{2{p3_bit_slice_38269_comb[13]}}, p3_bit_slice_38269_comb} - p2_sign_ext_36774;
  assign p3_smul_38383_comb = smul16b_16b_x_16b(p3_smul_38333_comb, p2_sub_37443);
  assign p3_sub_38384_comb = {{2{p3_bit_slice_38273_comb[13]}}, p3_bit_slice_38273_comb} - p2_sign_ext_36779;
  assign p3_smul_38387_comb = smul16b_16b_x_16b(p3_smul_38336_comb, p2_sub_37445);
  assign p3_sub_38388_comb = {{2{p3_bit_slice_38277_comb[13]}}, p3_bit_slice_38277_comb} - p2_sign_ext_36784;
  assign p3_smul_38391_comb = smul16b_16b_x_16b(p3_smul_38339_comb, p2_sub_37447);
  assign p3_sub_38392_comb = {{2{p3_bit_slice_38281_comb[13]}}, p3_bit_slice_38281_comb} - p2_sign_ext_36789;
  assign p3_smul_38395_comb = smul16b_16b_x_16b(p3_smul_38342_comb, p2_sub_37449);
  assign p3_sub_38396_comb = {{2{p3_bit_slice_38285_comb[13]}}, p3_bit_slice_38285_comb} - p2_sign_ext_36794;
  assign p3_smul_38399_comb = smul16b_16b_x_16b(p3_smul_38345_comb, p2_sub_37451);
  assign p3_sub_38400_comb = {{2{p3_bit_slice_38289_comb[13]}}, p3_bit_slice_38289_comb} - p2_sign_ext_36799;
  assign p3_smul_38403_comb = smul16b_16b_x_16b(p3_smul_38348_comb, p2_sub_37453);
  assign p3_sub_38404_comb = {{2{p3_bit_slice_38293_comb[13]}}, p3_bit_slice_38293_comb} - p2_sign_ext_36804;
  assign p3_add_38607_comb = p2_add_37551 + p2_add_37552;
  assign p3_add_38608_comb = p3_add_38559_comb + p3_add_38560_comb;
  assign p3_add_38609_comb = p3_smul_38127_comb + p3_smul_38183_comb;
  assign p3_add_38610_comb = p3_smul_38239_comb + p3_smul_38295_comb;
  assign p3_add_38611_comb = p2_add_37553 + p2_add_37554;
  assign p3_add_38612_comb = p3_add_38561_comb + p3_add_38562_comb;
  assign p3_add_38613_comb = p3_smul_38130_comb + p3_smul_38187_comb;
  assign p3_add_38614_comb = p3_smul_38242_comb + p3_smul_38299_comb;
  assign p3_add_38615_comb = p2_add_37555 + p2_add_37556;
  assign p3_add_38616_comb = p3_add_38563_comb + p3_add_38564_comb;
  assign p3_add_38617_comb = p3_smul_38133_comb + p3_smul_38191_comb;
  assign p3_add_38618_comb = p3_smul_38245_comb + p3_smul_38303_comb;
  assign p3_add_38619_comb = p2_add_37557 + p2_add_37558;
  assign p3_add_38620_comb = p3_add_38565_comb + p3_add_38566_comb;
  assign p3_add_38621_comb = p3_smul_38136_comb + p3_smul_38195_comb;
  assign p3_add_38622_comb = p3_smul_38248_comb + p3_smul_38307_comb;
  assign p3_add_38623_comb = p2_add_37559 + p2_add_37560;
  assign p3_add_38624_comb = p3_add_38567_comb + p3_add_38568_comb;
  assign p3_add_38625_comb = p3_smul_38139_comb + p3_smul_38199_comb;
  assign p3_add_38626_comb = p3_smul_38251_comb + p3_smul_38311_comb;
  assign p3_add_38627_comb = p2_add_37561 + p2_add_37562;
  assign p3_add_38628_comb = p3_add_38569_comb + p3_add_38570_comb;
  assign p3_add_38629_comb = p3_smul_38142_comb + p3_smul_38203_comb;
  assign p3_add_38630_comb = p3_smul_38254_comb + p3_smul_38315_comb;
  assign p3_add_38631_comb = p2_add_37563 + p2_add_37564;
  assign p3_add_38632_comb = p3_add_38571_comb + p3_add_38572_comb;
  assign p3_add_38633_comb = p3_smul_38145_comb + p3_smul_38207_comb;
  assign p3_add_38634_comb = p3_smul_38257_comb + p3_smul_38319_comb;
  assign p3_add_38635_comb = p2_add_37565 + p2_add_37566;
  assign p3_add_38636_comb = p3_add_38573_comb + p3_add_38574_comb;
  assign p3_add_38637_comb = p3_smul_38148_comb + p3_smul_38211_comb;
  assign p3_add_38638_comb = p3_smul_38260_comb + p3_smul_38323_comb;
  assign p3_add_38639_comb = p2_add_37567 + p3_add_38575_comb;
  assign p3_add_38640_comb = p3_add_38576_comb + p3_add_38577_comb;
  assign p3_add_38641_comb = p2_add_37568 + p3_add_38579_comb;
  assign p3_add_38642_comb = p3_add_38580_comb + p3_add_38581_comb;
  assign p3_add_38643_comb = p2_add_37569 + p3_add_38583_comb;
  assign p3_add_38644_comb = p3_add_38584_comb + p3_add_38585_comb;
  assign p3_add_38645_comb = p2_add_37570 + p3_add_38587_comb;
  assign p3_add_38646_comb = p3_add_38588_comb + p3_add_38589_comb;
  assign p3_add_38647_comb = p2_add_37571 + p3_add_38591_comb;
  assign p3_add_38648_comb = p3_add_38592_comb + p3_add_38593_comb;
  assign p3_add_38649_comb = p2_add_37572 + p3_add_38595_comb;
  assign p3_add_38650_comb = p3_add_38596_comb + p3_add_38597_comb;
  assign p3_add_38651_comb = p2_add_37573 + p3_add_38599_comb;
  assign p3_add_38652_comb = p3_add_38600_comb + p3_add_38601_comb;
  assign p3_add_38653_comb = p2_add_37574 + p3_add_38603_comb;
  assign p3_add_38654_comb = p3_add_38604_comb + p3_add_38605_comb;
  assign p3_smul_38407_comb = smul16b_16b_x_16b(p3_smul_38351_comb, p2_sub_37455);
  assign p3_sub_38408_comb = {{2{p3_bit_slice_38297_comb[13]}}, p3_bit_slice_38297_comb} - p2_sign_ext_36809;
  assign p3_smul_38411_comb = smul16b_16b_x_16b(p3_smul_38354_comb, p2_sub_37457);
  assign p3_sub_38412_comb = {{2{p3_bit_slice_38301_comb[13]}}, p3_bit_slice_38301_comb} - p2_sign_ext_36814;
  assign p3_smul_38415_comb = smul16b_16b_x_16b(p3_smul_38357_comb, p2_sub_37459);
  assign p3_sub_38416_comb = {{2{p3_bit_slice_38305_comb[13]}}, p3_bit_slice_38305_comb} - p2_sign_ext_36819;
  assign p3_smul_38419_comb = smul16b_16b_x_16b(p3_smul_38360_comb, p2_sub_37461);
  assign p3_sub_38420_comb = {{2{p3_bit_slice_38309_comb[13]}}, p3_bit_slice_38309_comb} - p2_sign_ext_36824;
  assign p3_smul_38423_comb = smul16b_16b_x_16b(p3_smul_38363_comb, p2_sub_37463);
  assign p3_sub_38424_comb = {{2{p3_bit_slice_38313_comb[13]}}, p3_bit_slice_38313_comb} - p2_sign_ext_36829;
  assign p3_smul_38427_comb = smul16b_16b_x_16b(p3_smul_38366_comb, p2_sub_37465);
  assign p3_sub_38428_comb = {{2{p3_bit_slice_38317_comb[13]}}, p3_bit_slice_38317_comb} - p2_sign_ext_36834;
  assign p3_smul_38431_comb = smul16b_16b_x_16b(p3_smul_38369_comb, p2_sub_37467);
  assign p3_sub_38432_comb = {{2{p3_bit_slice_38321_comb[13]}}, p3_bit_slice_38321_comb} - p2_sign_ext_36839;
  assign p3_smul_38435_comb = smul16b_16b_x_16b(p3_smul_38372_comb, p2_sub_37469);
  assign p3_sub_38436_comb = {{2{p3_bit_slice_38325_comb[13]}}, p3_bit_slice_38325_comb} - p2_sign_ext_36844;
  assign p3_smul_38439_comb = smul16b_16b_x_16b(p3_smul_38375_comb, p3_sub_38376_comb);
  assign p3_smul_38442_comb = smul16b_16b_x_16b(p3_smul_38379_comb, p3_sub_38380_comb);
  assign p3_smul_38445_comb = smul16b_16b_x_16b(p3_smul_38383_comb, p3_sub_38384_comb);
  assign p3_smul_38448_comb = smul16b_16b_x_16b(p3_smul_38387_comb, p3_sub_38388_comb);
  assign p3_smul_38451_comb = smul16b_16b_x_16b(p3_smul_38391_comb, p3_sub_38392_comb);
  assign p3_smul_38454_comb = smul16b_16b_x_16b(p3_smul_38395_comb, p3_sub_38396_comb);
  assign p3_smul_38457_comb = smul16b_16b_x_16b(p3_smul_38399_comb, p3_sub_38400_comb);
  assign p3_smul_38460_comb = smul16b_16b_x_16b(p3_smul_38403_comb, p3_sub_38404_comb);
  assign p3_sub_38479_comb = {{3{p3_bit_slice_38377_comb[12]}}, p3_bit_slice_38377_comb} - p2_sign_ext_36769;
  assign p3_sub_38481_comb = {{3{p3_bit_slice_38381_comb[12]}}, p3_bit_slice_38381_comb} - p2_sign_ext_36774;
  assign p3_sub_38483_comb = {{3{p3_bit_slice_38385_comb[12]}}, p3_bit_slice_38385_comb} - p2_sign_ext_36779;
  assign p3_sub_38485_comb = {{3{p3_bit_slice_38389_comb[12]}}, p3_bit_slice_38389_comb} - p2_sign_ext_36784;
  assign p3_sub_38487_comb = {{3{p3_bit_slice_38393_comb[12]}}, p3_bit_slice_38393_comb} - p2_sign_ext_36789;
  assign p3_sub_38489_comb = {{3{p3_bit_slice_38397_comb[12]}}, p3_bit_slice_38397_comb} - p2_sign_ext_36794;
  assign p3_sub_38491_comb = {{3{p3_bit_slice_38401_comb[12]}}, p3_bit_slice_38401_comb} - p2_sign_ext_36799;
  assign p3_sub_38493_comb = {{3{p3_bit_slice_38405_comb[12]}}, p3_bit_slice_38405_comb} - p2_sign_ext_36804;
  assign p3_sub_38495_comb = {{3{p3_bit_slice_38409_comb[12]}}, p3_bit_slice_38409_comb} - p2_sign_ext_36809;
  assign p3_sub_38497_comb = {{3{p3_bit_slice_38413_comb[12]}}, p3_bit_slice_38413_comb} - p2_sign_ext_36814;
  assign p3_sub_38499_comb = {{3{p3_bit_slice_38417_comb[12]}}, p3_bit_slice_38417_comb} - p2_sign_ext_36819;
  assign p3_sub_38501_comb = {{3{p3_bit_slice_38421_comb[12]}}, p3_bit_slice_38421_comb} - p2_sign_ext_36824;
  assign p3_sub_38503_comb = {{3{p3_bit_slice_38425_comb[12]}}, p3_bit_slice_38425_comb} - p2_sign_ext_36829;
  assign p3_sub_38505_comb = {{3{p3_bit_slice_38429_comb[12]}}, p3_bit_slice_38429_comb} - p2_sign_ext_36834;
  assign p3_sub_38507_comb = {{3{p3_bit_slice_38433_comb[12]}}, p3_bit_slice_38433_comb} - p2_sign_ext_36839;
  assign p3_sub_38509_comb = {{3{p3_bit_slice_38437_comb[12]}}, p3_bit_slice_38437_comb} - p2_sign_ext_36844;
  assign p3_sub_38527_comb = {{3{p3_bit_slice_38480_comb[12]}}, p3_bit_slice_38480_comb} - p2_sign_ext_36769;
  assign p3_sub_38528_comb = {{3{p3_bit_slice_38482_comb[12]}}, p3_bit_slice_38482_comb} - p2_sign_ext_36774;
  assign p3_sub_38529_comb = {{3{p3_bit_slice_38484_comb[12]}}, p3_bit_slice_38484_comb} - p2_sign_ext_36779;
  assign p3_sub_38530_comb = {{3{p3_bit_slice_38486_comb[12]}}, p3_bit_slice_38486_comb} - p2_sign_ext_36784;
  assign p3_sub_38531_comb = {{3{p3_bit_slice_38488_comb[12]}}, p3_bit_slice_38488_comb} - p2_sign_ext_36789;
  assign p3_sub_38532_comb = {{3{p3_bit_slice_38490_comb[12]}}, p3_bit_slice_38490_comb} - p2_sign_ext_36794;
  assign p3_sub_38533_comb = {{3{p3_bit_slice_38492_comb[12]}}, p3_bit_slice_38492_comb} - p2_sign_ext_36799;
  assign p3_sub_38534_comb = {{3{p3_bit_slice_38494_comb[12]}}, p3_bit_slice_38494_comb} - p2_sign_ext_36804;
  assign p3_sub_38535_comb = {{3{p3_bit_slice_38496_comb[12]}}, p3_bit_slice_38496_comb} - p2_sign_ext_36809;
  assign p3_sub_38536_comb = {{3{p3_bit_slice_38498_comb[12]}}, p3_bit_slice_38498_comb} - p2_sign_ext_36814;
  assign p3_sub_38537_comb = {{3{p3_bit_slice_38500_comb[12]}}, p3_bit_slice_38500_comb} - p2_sign_ext_36819;
  assign p3_sub_38538_comb = {{3{p3_bit_slice_38502_comb[12]}}, p3_bit_slice_38502_comb} - p2_sign_ext_36824;
  assign p3_sub_38539_comb = {{3{p3_bit_slice_38504_comb[12]}}, p3_bit_slice_38504_comb} - p2_sign_ext_36829;
  assign p3_sub_38540_comb = {{3{p3_bit_slice_38506_comb[12]}}, p3_bit_slice_38506_comb} - p2_sign_ext_36834;
  assign p3_sub_38541_comb = {{3{p3_bit_slice_38508_comb[12]}}, p3_bit_slice_38508_comb} - p2_sign_ext_36839;
  assign p3_sub_38542_comb = {{3{p3_bit_slice_38510_comb[12]}}, p3_bit_slice_38510_comb} - p2_sign_ext_36844;
  assign p3_add_38578_comb = p3_smul_38327_comb + p3_smul_38375_comb;
  assign p3_add_38582_comb = p3_smul_38330_comb + p3_smul_38379_comb;
  assign p3_add_38586_comb = p3_smul_38333_comb + p3_smul_38383_comb;
  assign p3_add_38590_comb = p3_smul_38336_comb + p3_smul_38387_comb;
  assign p3_add_38594_comb = p3_smul_38339_comb + p3_smul_38391_comb;
  assign p3_add_38598_comb = p3_smul_38342_comb + p3_smul_38395_comb;
  assign p3_add_38602_comb = p3_smul_38345_comb + p3_smul_38399_comb;
  assign p3_add_38606_comb = p3_smul_38348_comb + p3_smul_38403_comb;
  assign p3_add_38655_comb = p3_add_38607_comb + p3_add_38608_comb;
  assign p3_add_38656_comb = p3_add_38609_comb + p3_add_38610_comb;
  assign p3_add_38657_comb = p3_add_38611_comb + p3_add_38612_comb;
  assign p3_add_38658_comb = p3_add_38613_comb + p3_add_38614_comb;
  assign p3_add_38659_comb = p3_add_38615_comb + p3_add_38616_comb;
  assign p3_add_38660_comb = p3_add_38617_comb + p3_add_38618_comb;
  assign p3_add_38661_comb = p3_add_38619_comb + p3_add_38620_comb;
  assign p3_add_38662_comb = p3_add_38621_comb + p3_add_38622_comb;
  assign p3_add_38663_comb = p3_add_38623_comb + p3_add_38624_comb;
  assign p3_add_38664_comb = p3_add_38625_comb + p3_add_38626_comb;
  assign p3_add_38665_comb = p3_add_38627_comb + p3_add_38628_comb;
  assign p3_add_38666_comb = p3_add_38629_comb + p3_add_38630_comb;
  assign p3_add_38667_comb = p3_add_38631_comb + p3_add_38632_comb;
  assign p3_add_38668_comb = p3_add_38633_comb + p3_add_38634_comb;
  assign p3_add_38669_comb = p3_add_38635_comb + p3_add_38636_comb;
  assign p3_add_38670_comb = p3_add_38637_comb + p3_add_38638_comb;
  assign p3_add_38671_comb = p3_add_38639_comb + p3_add_38640_comb;
  assign p3_add_38672_comb = p3_add_38641_comb + p3_add_38642_comb;
  assign p3_add_38673_comb = p3_add_38643_comb + p3_add_38644_comb;
  assign p3_add_38674_comb = p3_add_38645_comb + p3_add_38646_comb;
  assign p3_add_38675_comb = p3_add_38647_comb + p3_add_38648_comb;
  assign p3_add_38676_comb = p3_add_38649_comb + p3_add_38650_comb;
  assign p3_add_38677_comb = p3_add_38651_comb + p3_add_38652_comb;
  assign p3_add_38678_comb = p3_add_38653_comb + p3_add_38654_comb;

  // Registers for pipe stage 3:
  reg [15:0] p3_smul_38351;
  reg [15:0] p3_smul_38354;
  reg [15:0] p3_smul_38357;
  reg [15:0] p3_smul_38360;
  reg [15:0] p3_smul_38363;
  reg [15:0] p3_smul_38366;
  reg [15:0] p3_smul_38369;
  reg [15:0] p3_smul_38372;
  reg [15:0] p3_smul_38407;
  reg [15:0] p3_sub_38408;
  reg [15:0] p3_smul_38411;
  reg [15:0] p3_sub_38412;
  reg [15:0] p3_smul_38415;
  reg [15:0] p3_sub_38416;
  reg [15:0] p3_smul_38419;
  reg [15:0] p3_sub_38420;
  reg [15:0] p3_smul_38423;
  reg [15:0] p3_sub_38424;
  reg [15:0] p3_smul_38427;
  reg [15:0] p3_sub_38428;
  reg [15:0] p3_smul_38431;
  reg [15:0] p3_sub_38432;
  reg [15:0] p3_smul_38435;
  reg [15:0] p3_sub_38436;
  reg [15:0] p3_smul_38439;
  reg [15:0] p3_bit_slice_37487;
  reg [15:0] p3_smul_38442;
  reg [15:0] p3_bit_slice_37488;
  reg [15:0] p3_smul_38445;
  reg [15:0] p3_bit_slice_37489;
  reg [15:0] p3_smul_38448;
  reg [15:0] p3_bit_slice_37490;
  reg [15:0] p3_smul_38451;
  reg [15:0] p3_bit_slice_37491;
  reg [15:0] p3_smul_38454;
  reg [15:0] p3_bit_slice_37492;
  reg [15:0] p3_smul_38457;
  reg [15:0] p3_bit_slice_37493;
  reg [15:0] p3_smul_38460;
  reg [15:0] p3_bit_slice_37494;
  reg [15:0] p3_bit_slice_37495;
  reg [15:0] p3_bit_slice_37496;
  reg [15:0] p3_bit_slice_37497;
  reg [15:0] p3_bit_slice_37498;
  reg [15:0] p3_bit_slice_37499;
  reg [15:0] p3_bit_slice_37500;
  reg [15:0] p3_bit_slice_37501;
  reg [15:0] p3_bit_slice_37502;
  reg [15:0] p3_sub_38479;
  reg [15:0] p3_sub_38481;
  reg [15:0] p3_sub_38483;
  reg [15:0] p3_sub_38485;
  reg [15:0] p3_sub_38487;
  reg [15:0] p3_sub_38489;
  reg [15:0] p3_sub_38491;
  reg [15:0] p3_sub_38493;
  reg [15:0] p3_sub_38495;
  reg [15:0] p3_sub_38497;
  reg [15:0] p3_sub_38499;
  reg [15:0] p3_sub_38501;
  reg [15:0] p3_sub_38503;
  reg [15:0] p3_sub_38505;
  reg [15:0] p3_sub_38507;
  reg [15:0] p3_sub_38509;
  reg [15:0] p3_sub_37519;
  reg [15:0] p3_sub_37520;
  reg [15:0] p3_sub_37521;
  reg [15:0] p3_sub_37522;
  reg [15:0] p3_sub_37523;
  reg [15:0] p3_sub_37524;
  reg [15:0] p3_sub_37525;
  reg [15:0] p3_sub_37526;
  reg [15:0] p3_sub_37527;
  reg [15:0] p3_sub_37528;
  reg [15:0] p3_sub_37529;
  reg [15:0] p3_sub_37530;
  reg [15:0] p3_sub_37531;
  reg [15:0] p3_sub_37532;
  reg [15:0] p3_sub_37533;
  reg [15:0] p3_sub_37534;
  reg [15:0] p3_sub_38527;
  reg [15:0] p3_sub_38528;
  reg [15:0] p3_sub_38529;
  reg [15:0] p3_sub_38530;
  reg [15:0] p3_sub_38531;
  reg [15:0] p3_sub_38532;
  reg [15:0] p3_sub_38533;
  reg [15:0] p3_sub_38534;
  reg [15:0] p3_sub_38535;
  reg [15:0] p3_sub_38536;
  reg [15:0] p3_sub_38537;
  reg [15:0] p3_sub_38538;
  reg [15:0] p3_sub_38539;
  reg [15:0] p3_sub_38540;
  reg [15:0] p3_sub_38541;
  reg [15:0] p3_sub_38542;
  reg [15:0] p3_add_38578;
  reg [15:0] p3_add_38582;
  reg [15:0] p3_add_38586;
  reg [15:0] p3_add_38590;
  reg [15:0] p3_add_38594;
  reg [15:0] p3_add_38598;
  reg [15:0] p3_add_38602;
  reg [15:0] p3_add_38606;
  reg [15:0] p3_add_38655;
  reg [15:0] p3_add_38656;
  reg [15:0] p3_add_38657;
  reg [15:0] p3_add_38658;
  reg [15:0] p3_add_38659;
  reg [15:0] p3_add_38660;
  reg [15:0] p3_add_38661;
  reg [15:0] p3_add_38662;
  reg [15:0] p3_add_38663;
  reg [15:0] p3_add_38664;
  reg [15:0] p3_add_38665;
  reg [15:0] p3_add_38666;
  reg [15:0] p3_add_38667;
  reg [15:0] p3_add_38668;
  reg [15:0] p3_add_38669;
  reg [15:0] p3_add_38670;
  reg [15:0] p3_add_38671;
  reg [15:0] p3_add_38672;
  reg [15:0] p3_add_38673;
  reg [15:0] p3_add_38674;
  reg [15:0] p3_add_38675;
  reg [15:0] p3_add_38676;
  reg [15:0] p3_add_38677;
  reg [15:0] p3_add_38678;
  always_ff @ (posedge clk) begin
    p3_smul_38351 <= p3_smul_38351_comb;
    p3_smul_38354 <= p3_smul_38354_comb;
    p3_smul_38357 <= p3_smul_38357_comb;
    p3_smul_38360 <= p3_smul_38360_comb;
    p3_smul_38363 <= p3_smul_38363_comb;
    p3_smul_38366 <= p3_smul_38366_comb;
    p3_smul_38369 <= p3_smul_38369_comb;
    p3_smul_38372 <= p3_smul_38372_comb;
    p3_smul_38407 <= p3_smul_38407_comb;
    p3_sub_38408 <= p3_sub_38408_comb;
    p3_smul_38411 <= p3_smul_38411_comb;
    p3_sub_38412 <= p3_sub_38412_comb;
    p3_smul_38415 <= p3_smul_38415_comb;
    p3_sub_38416 <= p3_sub_38416_comb;
    p3_smul_38419 <= p3_smul_38419_comb;
    p3_sub_38420 <= p3_sub_38420_comb;
    p3_smul_38423 <= p3_smul_38423_comb;
    p3_sub_38424 <= p3_sub_38424_comb;
    p3_smul_38427 <= p3_smul_38427_comb;
    p3_sub_38428 <= p3_sub_38428_comb;
    p3_smul_38431 <= p3_smul_38431_comb;
    p3_sub_38432 <= p3_sub_38432_comb;
    p3_smul_38435 <= p3_smul_38435_comb;
    p3_sub_38436 <= p3_sub_38436_comb;
    p3_smul_38439 <= p3_smul_38439_comb;
    p3_bit_slice_37487 <= p2_bit_slice_37487;
    p3_smul_38442 <= p3_smul_38442_comb;
    p3_bit_slice_37488 <= p2_bit_slice_37488;
    p3_smul_38445 <= p3_smul_38445_comb;
    p3_bit_slice_37489 <= p2_bit_slice_37489;
    p3_smul_38448 <= p3_smul_38448_comb;
    p3_bit_slice_37490 <= p2_bit_slice_37490;
    p3_smul_38451 <= p3_smul_38451_comb;
    p3_bit_slice_37491 <= p2_bit_slice_37491;
    p3_smul_38454 <= p3_smul_38454_comb;
    p3_bit_slice_37492 <= p2_bit_slice_37492;
    p3_smul_38457 <= p3_smul_38457_comb;
    p3_bit_slice_37493 <= p2_bit_slice_37493;
    p3_smul_38460 <= p3_smul_38460_comb;
    p3_bit_slice_37494 <= p2_bit_slice_37494;
    p3_bit_slice_37495 <= p2_bit_slice_37495;
    p3_bit_slice_37496 <= p2_bit_slice_37496;
    p3_bit_slice_37497 <= p2_bit_slice_37497;
    p3_bit_slice_37498 <= p2_bit_slice_37498;
    p3_bit_slice_37499 <= p2_bit_slice_37499;
    p3_bit_slice_37500 <= p2_bit_slice_37500;
    p3_bit_slice_37501 <= p2_bit_slice_37501;
    p3_bit_slice_37502 <= p2_bit_slice_37502;
    p3_sub_38479 <= p3_sub_38479_comb;
    p3_sub_38481 <= p3_sub_38481_comb;
    p3_sub_38483 <= p3_sub_38483_comb;
    p3_sub_38485 <= p3_sub_38485_comb;
    p3_sub_38487 <= p3_sub_38487_comb;
    p3_sub_38489 <= p3_sub_38489_comb;
    p3_sub_38491 <= p3_sub_38491_comb;
    p3_sub_38493 <= p3_sub_38493_comb;
    p3_sub_38495 <= p3_sub_38495_comb;
    p3_sub_38497 <= p3_sub_38497_comb;
    p3_sub_38499 <= p3_sub_38499_comb;
    p3_sub_38501 <= p3_sub_38501_comb;
    p3_sub_38503 <= p3_sub_38503_comb;
    p3_sub_38505 <= p3_sub_38505_comb;
    p3_sub_38507 <= p3_sub_38507_comb;
    p3_sub_38509 <= p3_sub_38509_comb;
    p3_sub_37519 <= p2_sub_37519;
    p3_sub_37520 <= p2_sub_37520;
    p3_sub_37521 <= p2_sub_37521;
    p3_sub_37522 <= p2_sub_37522;
    p3_sub_37523 <= p2_sub_37523;
    p3_sub_37524 <= p2_sub_37524;
    p3_sub_37525 <= p2_sub_37525;
    p3_sub_37526 <= p2_sub_37526;
    p3_sub_37527 <= p2_sub_37527;
    p3_sub_37528 <= p2_sub_37528;
    p3_sub_37529 <= p2_sub_37529;
    p3_sub_37530 <= p2_sub_37530;
    p3_sub_37531 <= p2_sub_37531;
    p3_sub_37532 <= p2_sub_37532;
    p3_sub_37533 <= p2_sub_37533;
    p3_sub_37534 <= p2_sub_37534;
    p3_sub_38527 <= p3_sub_38527_comb;
    p3_sub_38528 <= p3_sub_38528_comb;
    p3_sub_38529 <= p3_sub_38529_comb;
    p3_sub_38530 <= p3_sub_38530_comb;
    p3_sub_38531 <= p3_sub_38531_comb;
    p3_sub_38532 <= p3_sub_38532_comb;
    p3_sub_38533 <= p3_sub_38533_comb;
    p3_sub_38534 <= p3_sub_38534_comb;
    p3_sub_38535 <= p3_sub_38535_comb;
    p3_sub_38536 <= p3_sub_38536_comb;
    p3_sub_38537 <= p3_sub_38537_comb;
    p3_sub_38538 <= p3_sub_38538_comb;
    p3_sub_38539 <= p3_sub_38539_comb;
    p3_sub_38540 <= p3_sub_38540_comb;
    p3_sub_38541 <= p3_sub_38541_comb;
    p3_sub_38542 <= p3_sub_38542_comb;
    p3_add_38578 <= p3_add_38578_comb;
    p3_add_38582 <= p3_add_38582_comb;
    p3_add_38586 <= p3_add_38586_comb;
    p3_add_38590 <= p3_add_38590_comb;
    p3_add_38594 <= p3_add_38594_comb;
    p3_add_38598 <= p3_add_38598_comb;
    p3_add_38602 <= p3_add_38602_comb;
    p3_add_38606 <= p3_add_38606_comb;
    p3_add_38655 <= p3_add_38655_comb;
    p3_add_38656 <= p3_add_38656_comb;
    p3_add_38657 <= p3_add_38657_comb;
    p3_add_38658 <= p3_add_38658_comb;
    p3_add_38659 <= p3_add_38659_comb;
    p3_add_38660 <= p3_add_38660_comb;
    p3_add_38661 <= p3_add_38661_comb;
    p3_add_38662 <= p3_add_38662_comb;
    p3_add_38663 <= p3_add_38663_comb;
    p3_add_38664 <= p3_add_38664_comb;
    p3_add_38665 <= p3_add_38665_comb;
    p3_add_38666 <= p3_add_38666_comb;
    p3_add_38667 <= p3_add_38667_comb;
    p3_add_38668 <= p3_add_38668_comb;
    p3_add_38669 <= p3_add_38669_comb;
    p3_add_38670 <= p3_add_38670_comb;
    p3_add_38671 <= p3_add_38671_comb;
    p3_add_38672 <= p3_add_38672_comb;
    p3_add_38673 <= p3_add_38673_comb;
    p3_add_38674 <= p3_add_38674_comb;
    p3_add_38675 <= p3_add_38675_comb;
    p3_add_38676 <= p3_add_38676_comb;
    p3_add_38677 <= p3_add_38677_comb;
    p3_add_38678 <= p3_add_38678_comb;
  end

  // ===== Pipe stage 4:
  wire [15:0] p4_smul_38935_comb;
  wire [15:0] p4_smul_38936_comb;
  wire [15:0] p4_smul_38937_comb;
  wire [15:0] p4_smul_38938_comb;
  wire [15:0] p4_smul_38939_comb;
  wire [15:0] p4_smul_38940_comb;
  wire [15:0] p4_smul_38941_comb;
  wire [15:0] p4_smul_38942_comb;
  wire [15:0] p4_smul_38943_comb;
  wire [15:0] p4_smul_38944_comb;
  wire [15:0] p4_smul_38945_comb;
  wire [15:0] p4_smul_38946_comb;
  wire [15:0] p4_smul_38947_comb;
  wire [15:0] p4_smul_38948_comb;
  wire [15:0] p4_smul_38949_comb;
  wire [15:0] p4_smul_38950_comb;
  wire [15:0] p4_smul_38951_comb;
  wire [15:0] p4_smul_38952_comb;
  wire [15:0] p4_smul_38953_comb;
  wire [15:0] p4_smul_38954_comb;
  wire [15:0] p4_smul_38955_comb;
  wire [15:0] p4_smul_38956_comb;
  wire [15:0] p4_smul_38957_comb;
  wire [15:0] p4_smul_38958_comb;
  wire [15:0] p4_smul_38959_comb;
  wire [15:0] p4_smul_38960_comb;
  wire [15:0] p4_smul_38961_comb;
  wire [15:0] p4_smul_38962_comb;
  wire [15:0] p4_smul_38963_comb;
  wire [15:0] p4_smul_38964_comb;
  wire [15:0] p4_smul_38965_comb;
  wire [15:0] p4_smul_38966_comb;
  wire [15:0] p4_smul_38967_comb;
  wire [15:0] p4_smul_38968_comb;
  wire [15:0] p4_smul_38969_comb;
  wire [15:0] p4_smul_38970_comb;
  wire [15:0] p4_smul_38971_comb;
  wire [15:0] p4_smul_38972_comb;
  wire [15:0] p4_smul_38973_comb;
  wire [15:0] p4_smul_38974_comb;
  wire [15:0] p4_smul_38975_comb;
  wire [15:0] p4_smul_38976_comb;
  wire [15:0] p4_smul_38977_comb;
  wire [15:0] p4_smul_38978_comb;
  wire [15:0] p4_smul_38979_comb;
  wire [15:0] p4_smul_38980_comb;
  wire [15:0] p4_smul_38981_comb;
  wire [15:0] p4_smul_38982_comb;
  wire [15:0] p4_smul_38983_comb;
  wire [15:0] p4_smul_38984_comb;
  wire [15:0] p4_smul_38985_comb;
  wire [15:0] p4_smul_38986_comb;
  wire [15:0] p4_smul_38987_comb;
  wire [15:0] p4_smul_38988_comb;
  wire [15:0] p4_smul_38989_comb;
  wire [15:0] p4_smul_38990_comb;
  wire [15:0] p4_smul_38991_comb;
  wire [15:0] p4_smul_38993_comb;
  wire [15:0] p4_smul_38995_comb;
  wire [15:0] p4_smul_38997_comb;
  wire [15:0] p4_smul_38999_comb;
  wire [15:0] p4_smul_39001_comb;
  wire [15:0] p4_smul_39003_comb;
  wire [15:0] p4_smul_39005_comb;
  wire [15:0] p4_smul_39007_comb;
  wire [15:0] p4_smul_39009_comb;
  wire [15:0] p4_smul_39011_comb;
  wire [15:0] p4_smul_39013_comb;
  wire [15:0] p4_smul_39015_comb;
  wire [15:0] p4_smul_39017_comb;
  wire [15:0] p4_smul_39019_comb;
  wire [15:0] p4_smul_39021_comb;
  wire [15:0] p4_add_39023_comb;
  wire [15:0] p4_add_39024_comb;
  wire [15:0] p4_add_39025_comb;
  wire [15:0] p4_add_39026_comb;
  wire [15:0] p4_add_39027_comb;
  wire [15:0] p4_add_39028_comb;
  wire [15:0] p4_add_39029_comb;
  wire [15:0] p4_add_39030_comb;
  wire [15:0] p4_add_39031_comb;
  wire [15:0] p4_add_39032_comb;
  wire [15:0] p4_add_39033_comb;
  wire [15:0] p4_add_39034_comb;
  wire [15:0] p4_add_39035_comb;
  wire [15:0] p4_add_39036_comb;
  wire [15:0] p4_add_39037_comb;
  wire [15:0] p4_add_39038_comb;
  wire [15:0] p4_add_39039_comb;
  wire [15:0] p4_add_39040_comb;
  wire [15:0] p4_add_39041_comb;
  wire [15:0] p4_add_39042_comb;
  wire [15:0] p4_add_39043_comb;
  wire [15:0] p4_add_39044_comb;
  wire [15:0] p4_add_39045_comb;
  wire [15:0] p4_add_39046_comb;
  wire [15:0] p4_add_39047_comb;
  wire [15:0] p4_add_39048_comb;
  wire [15:0] p4_add_39049_comb;
  wire [15:0] p4_add_39050_comb;
  wire [15:0] p4_add_39051_comb;
  wire [15:0] p4_add_39052_comb;
  wire [15:0] p4_add_39053_comb;
  wire [15:0] p4_add_39054_comb;
  wire [15:0] p4_add_39055_comb;
  wire [15:0] p4_add_39056_comb;
  wire [15:0] p4_add_39057_comb;
  wire [15:0] p4_add_39058_comb;
  wire [15:0] p4_add_39059_comb;
  wire [15:0] p4_add_39060_comb;
  wire [15:0] p4_add_39061_comb;
  wire [15:0] p4_add_39062_comb;
  wire [15:0] p4_add_39063_comb;
  wire [15:0] p4_add_39064_comb;
  wire [15:0] p4_add_39065_comb;
  wire [15:0] p4_add_39066_comb;
  wire [15:0] p4_add_39067_comb;
  wire [15:0] p4_add_39068_comb;
  wire [15:0] p4_add_39069_comb;
  wire [15:0] p4_add_39070_comb;
  wire [15:0] p4_add_39071_comb;
  wire [15:0] p4_add_39072_comb;
  wire [15:0] p4_add_39073_comb;
  wire [15:0] p4_add_39074_comb;
  wire [15:0] p4_add_39075_comb;
  wire [15:0] p4_add_39076_comb;
  wire [15:0] p4_add_39077_comb;
  wire [15:0] p4_add_39078_comb;
  wire [15:0] p4_add_39079_comb;
  wire [15:0] p4_add_39080_comb;
  wire [15:0] p4_add_39081_comb;
  wire [15:0] p4_add_39082_comb;
  wire [15:0] p4_add_39083_comb;
  wire [15:0] p4_add_39084_comb;
  wire [15:0] p4_add_39085_comb;
  wire [15:0] p4_add_39086_comb;
  wire [15:0] p4_add_39087_comb;
  wire [15:0] p4_add_39088_comb;
  wire [15:0] p4_add_39089_comb;
  wire [15:0] p4_add_39090_comb;
  wire [15:0] p4_add_39091_comb;
  wire [15:0] p4_add_39092_comb;
  wire [15:0] p4_add_39093_comb;
  wire [15:0] p4_add_39094_comb;
  wire [15:0] p4_add_39095_comb;
  wire [15:0] p4_add_39096_comb;
  wire [15:0] p4_add_39097_comb;
  wire [15:0] p4_add_39098_comb;
  wire [15:0] p4_add_39099_comb;
  wire [15:0] p4_add_39100_comb;
  wire [15:0] p4_add_39101_comb;
  wire [15:0] p4_add_39102_comb;
  wire [15:0] p4_add_39103_comb;
  wire [15:0] p4_add_39104_comb;
  wire [15:0] p4_add_39105_comb;
  wire [15:0] p4_add_39106_comb;
  wire [15:0] p4_add_39107_comb;
  wire [15:0] p4_add_39108_comb;
  wire [15:0] p4_add_39109_comb;
  wire [15:0] p4_add_39110_comb;
  wire [15:0] p4_add_39111_comb;
  wire [15:0] p4_add_39112_comb;
  wire [15:0] p4_add_39113_comb;
  wire [15:0] p4_add_39114_comb;
  wire [15:0] p4_add_39115_comb;
  wire [15:0] p4_add_39116_comb;
  wire [15:0] p4_add_39117_comb;
  wire [15:0] p4_add_39118_comb;
  wire [15:0] p4_add_39119_comb;
  wire [15:0] p4_add_39120_comb;
  wire [15:0] p4_add_39121_comb;
  wire [15:0] p4_add_39122_comb;
  wire [15:0] p4_add_39123_comb;
  wire [15:0] p4_add_39124_comb;
  wire [15:0] p4_add_39125_comb;
  wire [15:0] p4_add_39126_comb;
  wire [15:0] p4_add_39127_comb;
  wire [15:0] p4_add_39128_comb;
  wire [15:0] p4_add_39129_comb;
  wire [15:0] p4_add_39130_comb;
  wire [15:0] p4_add_39131_comb;
  wire [15:0] p4_add_39132_comb;
  wire [15:0] p4_add_39133_comb;
  wire [15:0] p4_add_39134_comb;
  wire [15:0] p4_add_39135_comb;
  wire [15:0] p4_add_39136_comb;
  wire [15:0] p4_add_39137_comb;
  wire [15:0] p4_add_39138_comb;
  wire [15:0] p4_add_39139_comb;
  wire [15:0] p4_add_39140_comb;
  wire [15:0] p4_add_39141_comb;
  wire [15:0] p4_add_39142_comb;
  wire [15:0] p4_add_39143_comb;
  wire [15:0] p4_add_39144_comb;
  wire [15:0] p4_add_39145_comb;
  wire [15:0] p4_add_39146_comb;
  wire [15:0] p4_add_39147_comb;
  wire [15:0] p4_add_39148_comb;
  wire [15:0] p4_add_39149_comb;
  wire [15:0] p4_add_39150_comb;
  assign p4_smul_38935_comb = smul16b_16b_x_16b(p3_smul_38407, p3_sub_38408);
  assign p4_smul_38936_comb = smul16b_16b_x_16b(p3_smul_38411, p3_sub_38412);
  assign p4_smul_38937_comb = smul16b_16b_x_16b(p3_smul_38415, p3_sub_38416);
  assign p4_smul_38938_comb = smul16b_16b_x_16b(p3_smul_38419, p3_sub_38420);
  assign p4_smul_38939_comb = smul16b_16b_x_16b(p3_smul_38423, p3_sub_38424);
  assign p4_smul_38940_comb = smul16b_16b_x_16b(p3_smul_38427, p3_sub_38428);
  assign p4_smul_38941_comb = smul16b_16b_x_16b(p3_smul_38431, p3_sub_38432);
  assign p4_smul_38942_comb = smul16b_16b_x_16b(p3_smul_38435, p3_sub_38436);
  assign p4_smul_38943_comb = smul16b_16b_x_16b(p3_smul_38439, p3_bit_slice_37487);
  assign p4_smul_38944_comb = smul16b_16b_x_16b(p3_smul_38442, p3_bit_slice_37488);
  assign p4_smul_38945_comb = smul16b_16b_x_16b(p3_smul_38445, p3_bit_slice_37489);
  assign p4_smul_38946_comb = smul16b_16b_x_16b(p3_smul_38448, p3_bit_slice_37490);
  assign p4_smul_38947_comb = smul16b_16b_x_16b(p3_smul_38451, p3_bit_slice_37491);
  assign p4_smul_38948_comb = smul16b_16b_x_16b(p3_smul_38454, p3_bit_slice_37492);
  assign p4_smul_38949_comb = smul16b_16b_x_16b(p3_smul_38457, p3_bit_slice_37493);
  assign p4_smul_38950_comb = smul16b_16b_x_16b(p3_smul_38460, p3_bit_slice_37494);
  assign p4_smul_38951_comb = smul16b_16b_x_16b(p4_smul_38935_comb, p3_bit_slice_37495);
  assign p4_smul_38952_comb = smul16b_16b_x_16b(p4_smul_38936_comb, p3_bit_slice_37496);
  assign p4_smul_38953_comb = smul16b_16b_x_16b(p4_smul_38937_comb, p3_bit_slice_37497);
  assign p4_smul_38954_comb = smul16b_16b_x_16b(p4_smul_38938_comb, p3_bit_slice_37498);
  assign p4_smul_38955_comb = smul16b_16b_x_16b(p4_smul_38939_comb, p3_bit_slice_37499);
  assign p4_smul_38956_comb = smul16b_16b_x_16b(p4_smul_38940_comb, p3_bit_slice_37500);
  assign p4_smul_38957_comb = smul16b_16b_x_16b(p4_smul_38941_comb, p3_bit_slice_37501);
  assign p4_smul_38958_comb = smul16b_16b_x_16b(p4_smul_38942_comb, p3_bit_slice_37502);
  assign p4_smul_38959_comb = smul16b_16b_x_16b(p4_smul_38943_comb, p3_sub_38479);
  assign p4_smul_38960_comb = smul16b_16b_x_16b(p4_smul_38944_comb, p3_sub_38481);
  assign p4_smul_38961_comb = smul16b_16b_x_16b(p4_smul_38945_comb, p3_sub_38483);
  assign p4_smul_38962_comb = smul16b_16b_x_16b(p4_smul_38946_comb, p3_sub_38485);
  assign p4_smul_38963_comb = smul16b_16b_x_16b(p4_smul_38947_comb, p3_sub_38487);
  assign p4_smul_38964_comb = smul16b_16b_x_16b(p4_smul_38948_comb, p3_sub_38489);
  assign p4_smul_38965_comb = smul16b_16b_x_16b(p4_smul_38949_comb, p3_sub_38491);
  assign p4_smul_38966_comb = smul16b_16b_x_16b(p4_smul_38950_comb, p3_sub_38493);
  assign p4_smul_38967_comb = smul16b_16b_x_16b(p4_smul_38951_comb, p3_sub_38495);
  assign p4_smul_38968_comb = smul16b_16b_x_16b(p4_smul_38952_comb, p3_sub_38497);
  assign p4_smul_38969_comb = smul16b_16b_x_16b(p4_smul_38953_comb, p3_sub_38499);
  assign p4_smul_38970_comb = smul16b_16b_x_16b(p4_smul_38954_comb, p3_sub_38501);
  assign p4_smul_38971_comb = smul16b_16b_x_16b(p4_smul_38955_comb, p3_sub_38503);
  assign p4_smul_38972_comb = smul16b_16b_x_16b(p4_smul_38956_comb, p3_sub_38505);
  assign p4_smul_38973_comb = smul16b_16b_x_16b(p4_smul_38957_comb, p3_sub_38507);
  assign p4_smul_38974_comb = smul16b_16b_x_16b(p4_smul_38958_comb, p3_sub_38509);
  assign p4_smul_38975_comb = smul16b_16b_x_16b(p4_smul_38959_comb, p3_sub_37519);
  assign p4_smul_38976_comb = smul16b_16b_x_16b(p4_smul_38960_comb, p3_sub_37520);
  assign p4_smul_38977_comb = smul16b_16b_x_16b(p4_smul_38961_comb, p3_sub_37521);
  assign p4_smul_38978_comb = smul16b_16b_x_16b(p4_smul_38962_comb, p3_sub_37522);
  assign p4_smul_38979_comb = smul16b_16b_x_16b(p4_smul_38963_comb, p3_sub_37523);
  assign p4_smul_38980_comb = smul16b_16b_x_16b(p4_smul_38964_comb, p3_sub_37524);
  assign p4_smul_38981_comb = smul16b_16b_x_16b(p4_smul_38965_comb, p3_sub_37525);
  assign p4_smul_38982_comb = smul16b_16b_x_16b(p4_smul_38966_comb, p3_sub_37526);
  assign p4_smul_38983_comb = smul16b_16b_x_16b(p4_smul_38967_comb, p3_sub_37527);
  assign p4_smul_38984_comb = smul16b_16b_x_16b(p4_smul_38968_comb, p3_sub_37528);
  assign p4_smul_38985_comb = smul16b_16b_x_16b(p4_smul_38969_comb, p3_sub_37529);
  assign p4_smul_38986_comb = smul16b_16b_x_16b(p4_smul_38970_comb, p3_sub_37530);
  assign p4_smul_38987_comb = smul16b_16b_x_16b(p4_smul_38971_comb, p3_sub_37531);
  assign p4_smul_38988_comb = smul16b_16b_x_16b(p4_smul_38972_comb, p3_sub_37532);
  assign p4_smul_38989_comb = smul16b_16b_x_16b(p4_smul_38973_comb, p3_sub_37533);
  assign p4_smul_38990_comb = smul16b_16b_x_16b(p4_smul_38974_comb, p3_sub_37534);
  assign p4_smul_38991_comb = smul16b_16b_x_16b(p4_smul_38975_comb, p3_sub_38527);
  assign p4_smul_38993_comb = smul16b_16b_x_16b(p4_smul_38976_comb, p3_sub_38528);
  assign p4_smul_38995_comb = smul16b_16b_x_16b(p4_smul_38977_comb, p3_sub_38529);
  assign p4_smul_38997_comb = smul16b_16b_x_16b(p4_smul_38978_comb, p3_sub_38530);
  assign p4_smul_38999_comb = smul16b_16b_x_16b(p4_smul_38979_comb, p3_sub_38531);
  assign p4_smul_39001_comb = smul16b_16b_x_16b(p4_smul_38980_comb, p3_sub_38532);
  assign p4_smul_39003_comb = smul16b_16b_x_16b(p4_smul_38981_comb, p3_sub_38533);
  assign p4_smul_39005_comb = smul16b_16b_x_16b(p4_smul_38982_comb, p3_sub_38534);
  assign p4_smul_39007_comb = smul16b_16b_x_16b(p4_smul_38983_comb, p3_sub_38535);
  assign p4_smul_39009_comb = smul16b_16b_x_16b(p4_smul_38984_comb, p3_sub_38536);
  assign p4_smul_39011_comb = smul16b_16b_x_16b(p4_smul_38985_comb, p3_sub_38537);
  assign p4_smul_39013_comb = smul16b_16b_x_16b(p4_smul_38986_comb, p3_sub_38538);
  assign p4_smul_39015_comb = smul16b_16b_x_16b(p4_smul_38987_comb, p3_sub_38539);
  assign p4_smul_39017_comb = smul16b_16b_x_16b(p4_smul_38988_comb, p3_sub_38540);
  assign p4_smul_39019_comb = smul16b_16b_x_16b(p4_smul_38989_comb, p3_sub_38541);
  assign p4_smul_39021_comb = smul16b_16b_x_16b(p4_smul_38990_comb, p3_sub_38542);
  assign p4_add_39023_comb = p3_smul_38439 + p4_smul_38943_comb;
  assign p4_add_39024_comb = p4_smul_38959_comb + p4_smul_38975_comb;
  assign p4_add_39025_comb = p4_smul_38991_comb + 16'h0001;
  assign p4_add_39026_comb = p3_smul_38442 + p4_smul_38944_comb;
  assign p4_add_39027_comb = p4_smul_38960_comb + p4_smul_38976_comb;
  assign p4_add_39028_comb = p4_smul_38993_comb + 16'h0001;
  assign p4_add_39029_comb = p3_smul_38445 + p4_smul_38945_comb;
  assign p4_add_39030_comb = p4_smul_38961_comb + p4_smul_38977_comb;
  assign p4_add_39031_comb = p4_smul_38995_comb + 16'h0001;
  assign p4_add_39032_comb = p3_smul_38448 + p4_smul_38946_comb;
  assign p4_add_39033_comb = p4_smul_38962_comb + p4_smul_38978_comb;
  assign p4_add_39034_comb = p4_smul_38997_comb + 16'h0001;
  assign p4_add_39035_comb = p3_smul_38451 + p4_smul_38947_comb;
  assign p4_add_39036_comb = p4_smul_38963_comb + p4_smul_38979_comb;
  assign p4_add_39037_comb = p4_smul_38999_comb + 16'h0001;
  assign p4_add_39038_comb = p3_smul_38454 + p4_smul_38948_comb;
  assign p4_add_39039_comb = p4_smul_38964_comb + p4_smul_38980_comb;
  assign p4_add_39040_comb = p4_smul_39001_comb + 16'h0001;
  assign p4_add_39041_comb = p3_smul_38457 + p4_smul_38949_comb;
  assign p4_add_39042_comb = p4_smul_38965_comb + p4_smul_38981_comb;
  assign p4_add_39043_comb = p4_smul_39003_comb + 16'h0001;
  assign p4_add_39044_comb = p3_smul_38460 + p4_smul_38950_comb;
  assign p4_add_39045_comb = p4_smul_38966_comb + p4_smul_38982_comb;
  assign p4_add_39046_comb = p4_smul_39005_comb + 16'h0001;
  assign p4_add_39047_comb = p3_smul_38351 + p3_smul_38407;
  assign p4_add_39048_comb = p4_smul_38935_comb + p4_smul_38951_comb;
  assign p4_add_39049_comb = p4_smul_38967_comb + p4_smul_38983_comb;
  assign p4_add_39050_comb = p4_smul_39007_comb + 16'h0001;
  assign p4_add_39051_comb = p3_smul_38354 + p3_smul_38411;
  assign p4_add_39052_comb = p4_smul_38936_comb + p4_smul_38952_comb;
  assign p4_add_39053_comb = p4_smul_38968_comb + p4_smul_38984_comb;
  assign p4_add_39054_comb = p4_smul_39009_comb + 16'h0001;
  assign p4_add_39055_comb = p3_smul_38357 + p3_smul_38415;
  assign p4_add_39056_comb = p4_smul_38937_comb + p4_smul_38953_comb;
  assign p4_add_39057_comb = p4_smul_38969_comb + p4_smul_38985_comb;
  assign p4_add_39058_comb = p4_smul_39011_comb + 16'h0001;
  assign p4_add_39059_comb = p3_smul_38360 + p3_smul_38419;
  assign p4_add_39060_comb = p4_smul_38938_comb + p4_smul_38954_comb;
  assign p4_add_39061_comb = p4_smul_38970_comb + p4_smul_38986_comb;
  assign p4_add_39062_comb = p4_smul_39013_comb + 16'h0001;
  assign p4_add_39063_comb = p3_smul_38363 + p3_smul_38423;
  assign p4_add_39064_comb = p4_smul_38939_comb + p4_smul_38955_comb;
  assign p4_add_39065_comb = p4_smul_38971_comb + p4_smul_38987_comb;
  assign p4_add_39066_comb = p4_smul_39015_comb + 16'h0001;
  assign p4_add_39067_comb = p3_smul_38366 + p3_smul_38427;
  assign p4_add_39068_comb = p4_smul_38940_comb + p4_smul_38956_comb;
  assign p4_add_39069_comb = p4_smul_38972_comb + p4_smul_38988_comb;
  assign p4_add_39070_comb = p4_smul_39017_comb + 16'h0001;
  assign p4_add_39071_comb = p3_smul_38369 + p3_smul_38431;
  assign p4_add_39072_comb = p4_smul_38941_comb + p4_smul_38957_comb;
  assign p4_add_39073_comb = p4_smul_38973_comb + p4_smul_38989_comb;
  assign p4_add_39074_comb = p4_smul_39019_comb + 16'h0001;
  assign p4_add_39075_comb = p3_smul_38372 + p3_smul_38435;
  assign p4_add_39076_comb = p4_smul_38942_comb + p4_smul_38958_comb;
  assign p4_add_39077_comb = p4_smul_38974_comb + p4_smul_38990_comb;
  assign p4_add_39078_comb = p4_smul_39021_comb + 16'h0001;
  assign p4_add_39079_comb = p3_add_38578 + p4_add_39023_comb;
  assign p4_add_39080_comb = p4_add_39024_comb + p4_add_39025_comb;
  assign p4_add_39081_comb = p3_add_38582 + p4_add_39026_comb;
  assign p4_add_39082_comb = p4_add_39027_comb + p4_add_39028_comb;
  assign p4_add_39083_comb = p3_add_38586 + p4_add_39029_comb;
  assign p4_add_39084_comb = p4_add_39030_comb + p4_add_39031_comb;
  assign p4_add_39085_comb = p3_add_38590 + p4_add_39032_comb;
  assign p4_add_39086_comb = p4_add_39033_comb + p4_add_39034_comb;
  assign p4_add_39087_comb = p3_add_38594 + p4_add_39035_comb;
  assign p4_add_39088_comb = p4_add_39036_comb + p4_add_39037_comb;
  assign p4_add_39089_comb = p3_add_38598 + p4_add_39038_comb;
  assign p4_add_39090_comb = p4_add_39039_comb + p4_add_39040_comb;
  assign p4_add_39091_comb = p3_add_38602 + p4_add_39041_comb;
  assign p4_add_39092_comb = p4_add_39042_comb + p4_add_39043_comb;
  assign p4_add_39093_comb = p3_add_38606 + p4_add_39044_comb;
  assign p4_add_39094_comb = p4_add_39045_comb + p4_add_39046_comb;
  assign p4_add_39095_comb = p4_add_39047_comb + p4_add_39048_comb;
  assign p4_add_39096_comb = p4_add_39049_comb + p4_add_39050_comb;
  assign p4_add_39097_comb = p4_add_39051_comb + p4_add_39052_comb;
  assign p4_add_39098_comb = p4_add_39053_comb + p4_add_39054_comb;
  assign p4_add_39099_comb = p4_add_39055_comb + p4_add_39056_comb;
  assign p4_add_39100_comb = p4_add_39057_comb + p4_add_39058_comb;
  assign p4_add_39101_comb = p4_add_39059_comb + p4_add_39060_comb;
  assign p4_add_39102_comb = p4_add_39061_comb + p4_add_39062_comb;
  assign p4_add_39103_comb = p4_add_39063_comb + p4_add_39064_comb;
  assign p4_add_39104_comb = p4_add_39065_comb + p4_add_39066_comb;
  assign p4_add_39105_comb = p4_add_39067_comb + p4_add_39068_comb;
  assign p4_add_39106_comb = p4_add_39069_comb + p4_add_39070_comb;
  assign p4_add_39107_comb = p4_add_39071_comb + p4_add_39072_comb;
  assign p4_add_39108_comb = p4_add_39073_comb + p4_add_39074_comb;
  assign p4_add_39109_comb = p4_add_39075_comb + p4_add_39076_comb;
  assign p4_add_39110_comb = p4_add_39077_comb + p4_add_39078_comb;
  assign p4_add_39111_comb = p4_add_39079_comb + p4_add_39080_comb;
  assign p4_add_39112_comb = p4_add_39081_comb + p4_add_39082_comb;
  assign p4_add_39113_comb = p4_add_39083_comb + p4_add_39084_comb;
  assign p4_add_39114_comb = p4_add_39085_comb + p4_add_39086_comb;
  assign p4_add_39115_comb = p4_add_39087_comb + p4_add_39088_comb;
  assign p4_add_39116_comb = p4_add_39089_comb + p4_add_39090_comb;
  assign p4_add_39117_comb = p4_add_39091_comb + p4_add_39092_comb;
  assign p4_add_39118_comb = p4_add_39093_comb + p4_add_39094_comb;
  assign p4_add_39119_comb = p3_add_38655 + p3_add_38656;
  assign p4_add_39120_comb = p4_add_39095_comb + p4_add_39096_comb;
  assign p4_add_39121_comb = p3_add_38657 + p3_add_38658;
  assign p4_add_39122_comb = p4_add_39097_comb + p4_add_39098_comb;
  assign p4_add_39123_comb = p3_add_38659 + p3_add_38660;
  assign p4_add_39124_comb = p4_add_39099_comb + p4_add_39100_comb;
  assign p4_add_39125_comb = p3_add_38661 + p3_add_38662;
  assign p4_add_39126_comb = p4_add_39101_comb + p4_add_39102_comb;
  assign p4_add_39127_comb = p3_add_38663 + p3_add_38664;
  assign p4_add_39128_comb = p4_add_39103_comb + p4_add_39104_comb;
  assign p4_add_39129_comb = p3_add_38665 + p3_add_38666;
  assign p4_add_39130_comb = p4_add_39105_comb + p4_add_39106_comb;
  assign p4_add_39131_comb = p3_add_38667 + p3_add_38668;
  assign p4_add_39132_comb = p4_add_39107_comb + p4_add_39108_comb;
  assign p4_add_39133_comb = p3_add_38669 + p3_add_38670;
  assign p4_add_39134_comb = p4_add_39109_comb + p4_add_39110_comb;
  assign p4_add_39135_comb = p3_add_38671 + p4_add_39111_comb;
  assign p4_add_39136_comb = p3_add_38672 + p4_add_39112_comb;
  assign p4_add_39137_comb = p3_add_38673 + p4_add_39113_comb;
  assign p4_add_39138_comb = p3_add_38674 + p4_add_39114_comb;
  assign p4_add_39139_comb = p3_add_38675 + p4_add_39115_comb;
  assign p4_add_39140_comb = p3_add_38676 + p4_add_39116_comb;
  assign p4_add_39141_comb = p3_add_38677 + p4_add_39117_comb;
  assign p4_add_39142_comb = p3_add_38678 + p4_add_39118_comb;
  assign p4_add_39143_comb = p4_add_39119_comb + p4_add_39120_comb;
  assign p4_add_39144_comb = p4_add_39121_comb + p4_add_39122_comb;
  assign p4_add_39145_comb = p4_add_39123_comb + p4_add_39124_comb;
  assign p4_add_39146_comb = p4_add_39125_comb + p4_add_39126_comb;
  assign p4_add_39147_comb = p4_add_39127_comb + p4_add_39128_comb;
  assign p4_add_39148_comb = p4_add_39129_comb + p4_add_39130_comb;
  assign p4_add_39149_comb = p4_add_39131_comb + p4_add_39132_comb;
  assign p4_add_39150_comb = p4_add_39133_comb + p4_add_39134_comb;

  // Registers for pipe stage 4:
  reg [15:0] p4_add_39135;
  reg [15:0] p4_add_39136;
  reg [15:0] p4_add_39137;
  reg [15:0] p4_add_39138;
  reg [15:0] p4_add_39139;
  reg [15:0] p4_add_39140;
  reg [15:0] p4_add_39141;
  reg [15:0] p4_add_39142;
  reg [15:0] p4_add_39143;
  reg [15:0] p4_add_39144;
  reg [15:0] p4_add_39145;
  reg [15:0] p4_add_39146;
  reg [15:0] p4_add_39147;
  reg [15:0] p4_add_39148;
  reg [15:0] p4_add_39149;
  reg [15:0] p4_add_39150;
  always_ff @ (posedge clk) begin
    p4_add_39135 <= p4_add_39135_comb;
    p4_add_39136 <= p4_add_39136_comb;
    p4_add_39137 <= p4_add_39137_comb;
    p4_add_39138 <= p4_add_39138_comb;
    p4_add_39139 <= p4_add_39139_comb;
    p4_add_39140 <= p4_add_39140_comb;
    p4_add_39141 <= p4_add_39141_comb;
    p4_add_39142 <= p4_add_39142_comb;
    p4_add_39143 <= p4_add_39143_comb;
    p4_add_39144 <= p4_add_39144_comb;
    p4_add_39145 <= p4_add_39145_comb;
    p4_add_39146 <= p4_add_39146_comb;
    p4_add_39147 <= p4_add_39147_comb;
    p4_add_39148 <= p4_add_39148_comb;
    p4_add_39149 <= p4_add_39149_comb;
    p4_add_39150 <= p4_add_39150_comb;
  end

  // ===== Pipe stage 5:
  wire [31:0] p5_add_39216_comb;
  wire [31:0] p5_add_39218_comb;
  wire [31:0] p5_add_39220_comb;
  wire [31:0] p5_add_39222_comb;
  wire [31:0] p5_add_39224_comb;
  wire [31:0] p5_add_39226_comb;
  wire [31:0] p5_add_39228_comb;
  wire [31:0] p5_add_39230_comb;
  wire [31:0] p5_add_39232_comb;
  wire [31:0] p5_add_39234_comb;
  wire [31:0] p5_add_39236_comb;
  wire [31:0] p5_add_39238_comb;
  wire [31:0] p5_add_39240_comb;
  wire [31:0] p5_add_39242_comb;
  wire [31:0] p5_add_39244_comb;
  wire [31:0] p5_add_39246_comb;
  wire [31:0] p5_sdiv_39247_comb;
  wire [31:0] p5_sdiv_39248_comb;
  wire [31:0] p5_sdiv_39249_comb;
  wire [31:0] p5_sdiv_39250_comb;
  wire [31:0] p5_sdiv_39251_comb;
  wire [31:0] p5_sdiv_39252_comb;
  wire [31:0] p5_sdiv_39253_comb;
  wire [31:0] p5_sdiv_39254_comb;
  wire [31:0] p5_sdiv_39255_comb;
  wire [31:0] p5_sdiv_39256_comb;
  wire [31:0] p5_sdiv_39257_comb;
  wire [31:0] p5_sdiv_39258_comb;
  wire [31:0] p5_sdiv_39259_comb;
  wire [31:0] p5_sdiv_39260_comb;
  wire [31:0] p5_sdiv_39261_comb;
  wire [31:0] p5_sdiv_39262_comb;
  wire [15:0] p5_array_39279_comb[16];
  assign p5_add_39216_comb = {{16{p4_add_39135[15]}}, p4_add_39135} + 32'h0000_0001;
  assign p5_add_39218_comb = {{16{p4_add_39136[15]}}, p4_add_39136} + 32'h0000_0001;
  assign p5_add_39220_comb = {{16{p4_add_39137[15]}}, p4_add_39137} + 32'h0000_0001;
  assign p5_add_39222_comb = {{16{p4_add_39138[15]}}, p4_add_39138} + 32'h0000_0001;
  assign p5_add_39224_comb = {{16{p4_add_39139[15]}}, p4_add_39139} + 32'h0000_0001;
  assign p5_add_39226_comb = {{16{p4_add_39140[15]}}, p4_add_39140} + 32'h0000_0001;
  assign p5_add_39228_comb = {{16{p4_add_39141[15]}}, p4_add_39141} + 32'h0000_0001;
  assign p5_add_39230_comb = {{16{p4_add_39142[15]}}, p4_add_39142} + 32'h0000_0001;
  assign p5_add_39232_comb = {{16{p4_add_39143[15]}}, p4_add_39143} + 32'h0000_0001;
  assign p5_add_39234_comb = {{16{p4_add_39144[15]}}, p4_add_39144} + 32'h0000_0001;
  assign p5_add_39236_comb = {{16{p4_add_39145[15]}}, p4_add_39145} + 32'h0000_0001;
  assign p5_add_39238_comb = {{16{p4_add_39146[15]}}, p4_add_39146} + 32'h0000_0001;
  assign p5_add_39240_comb = {{16{p4_add_39147[15]}}, p4_add_39147} + 32'h0000_0001;
  assign p5_add_39242_comb = {{16{p4_add_39148[15]}}, p4_add_39148} + 32'h0000_0001;
  assign p5_add_39244_comb = {{16{p4_add_39149[15]}}, p4_add_39149} + 32'h0000_0001;
  assign p5_add_39246_comb = {{16{p4_add_39150[15]}}, p4_add_39150} + 32'h0000_0001;
  assign p5_sdiv_39247_comb = sdiv_32b(32'h0000_0001, p5_add_39216_comb);
  assign p5_sdiv_39248_comb = sdiv_32b(32'h0000_0001, p5_add_39218_comb);
  assign p5_sdiv_39249_comb = sdiv_32b(32'h0000_0001, p5_add_39220_comb);
  assign p5_sdiv_39250_comb = sdiv_32b(32'h0000_0001, p5_add_39222_comb);
  assign p5_sdiv_39251_comb = sdiv_32b(32'h0000_0001, p5_add_39224_comb);
  assign p5_sdiv_39252_comb = sdiv_32b(32'h0000_0001, p5_add_39226_comb);
  assign p5_sdiv_39253_comb = sdiv_32b(32'h0000_0001, p5_add_39228_comb);
  assign p5_sdiv_39254_comb = sdiv_32b(32'h0000_0001, p5_add_39230_comb);
  assign p5_sdiv_39255_comb = sdiv_32b(32'h0000_0001, p5_add_39232_comb);
  assign p5_sdiv_39256_comb = sdiv_32b(32'h0000_0001, p5_add_39234_comb);
  assign p5_sdiv_39257_comb = sdiv_32b(32'h0000_0001, p5_add_39236_comb);
  assign p5_sdiv_39258_comb = sdiv_32b(32'h0000_0001, p5_add_39238_comb);
  assign p5_sdiv_39259_comb = sdiv_32b(32'h0000_0001, p5_add_39240_comb);
  assign p5_sdiv_39260_comb = sdiv_32b(32'h0000_0001, p5_add_39242_comb);
  assign p5_sdiv_39261_comb = sdiv_32b(32'h0000_0001, p5_add_39244_comb);
  assign p5_sdiv_39262_comb = sdiv_32b(32'h0000_0001, p5_add_39246_comb);
  assign p5_array_39279_comb[0] = p5_sdiv_39247_comb[15:0];
  assign p5_array_39279_comb[1] = p5_sdiv_39248_comb[15:0];
  assign p5_array_39279_comb[2] = p5_sdiv_39249_comb[15:0];
  assign p5_array_39279_comb[3] = p5_sdiv_39250_comb[15:0];
  assign p5_array_39279_comb[4] = p5_sdiv_39251_comb[15:0];
  assign p5_array_39279_comb[5] = p5_sdiv_39252_comb[15:0];
  assign p5_array_39279_comb[6] = p5_sdiv_39253_comb[15:0];
  assign p5_array_39279_comb[7] = p5_sdiv_39254_comb[15:0];
  assign p5_array_39279_comb[8] = p5_sdiv_39255_comb[15:0];
  assign p5_array_39279_comb[9] = p5_sdiv_39256_comb[15:0];
  assign p5_array_39279_comb[10] = p5_sdiv_39257_comb[15:0];
  assign p5_array_39279_comb[11] = p5_sdiv_39258_comb[15:0];
  assign p5_array_39279_comb[12] = p5_sdiv_39259_comb[15:0];
  assign p5_array_39279_comb[13] = p5_sdiv_39260_comb[15:0];
  assign p5_array_39279_comb[14] = p5_sdiv_39261_comb[15:0];
  assign p5_array_39279_comb[15] = p5_sdiv_39262_comb[15:0];

  // Registers for pipe stage 5:
  reg [15:0] p5_array_39279[16];
  always_ff @ (posedge clk) begin
    p5_array_39279 <= p5_array_39279_comb;
  end
  assign out = {p5_array_39279[15], p5_array_39279[14], p5_array_39279[13], p5_array_39279[12], p5_array_39279[11], p5_array_39279[10], p5_array_39279[9], p5_array_39279[8], p5_array_39279[7], p5_array_39279[6], p5_array_39279[5], p5_array_39279[4], p5_array_39279[3], p5_array_39279[2], p5_array_39279[1], p5_array_39279[0]};
endmodule
